13087 24
18 1 2 3 4 5 6 7 8 9 10 10 11 10 12 13 14 15 16 
26 1 2 3 9 4 6 5 7 8 9 10 5 17 7 8 10 10 11 10 16 16 14 13 12 15 16 
37 1 2 3 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 5 17 7 8 10 10 10 10 10 10 11 10 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 19 9 
8 1 2 3 20 9 9 18 9 
8 1 2 3 9 9 9 9 19 
8 1 2 3 20 9 9 19 9 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 18 21 16 
43 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 14 13 12 15 16 
21 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 21 18 22 
11 1 2 20 3 20 9 9 9 9 18 9 
3 1 2 18 
40 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 22 22 16 22 22 16 22 22 22 16 16 14 15 12 13 16 
4 1 2 18 20 
35 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 11 10 16 22 22 22 5 17 7 8 22 22 11 22 14 13 12 15 16 
28 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 22 22 14 12 13 15 16 
21 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
13 1 2 3 20 4 5 6 7 8 9 17 19 10 
24 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 17 5 7 8 10 10 18 21 10 
17 1 2 3 9 4 6 5 7 8 9 11 10 14 12 15 13 16 
22 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 23 18 23 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 13 15 12 14 16 
4 1 2 18 20 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 18 9 
4 1 2 18 20 
5 1 2 3 18 9 
56 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 16 22 22 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 13 14 15 12 16 
23 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 19 17 10 
19 1 2 3 4 5 6 7 8 9 10 10 11 10 16 14 13 15 12 16 
22 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 16 14 12 15 13 16 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
8 1 2 3 9 9 9 18 9 
4 1 2 18 20 
25 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
28 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
6 1 2 3 20 18 9 
20 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 11 10 18 21 16 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 10 11 10 16 21 18 16 
11 1 2 20 20 3 20 9 9 9 18 9 
7 1 2 20 3 20 18 9 
3 1 2 18 
19 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
3 1 2 18 
7 1 2 3 9 9 19 9 
18 1 2 3 9 9 4 6 5 7 8 9 11 10 14 13 12 15 16 
14 1 2 3 4 6 5 7 8 9 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
14 1 2 3 20 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 21 18 16 
22 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 21 18 16 
3 1 2 18 
3 1 2 18 
36 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 11 10 16 16 22 17 5 7 8 22 22 22 22 11 22 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
17 1 2 3 20 9 9 4 6 5 7 8 9 10 10 17 19 10 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 14 15 13 12 16 
6 1 2 23 23 18 23 
10 1 2 3 20 9 9 9 9 19 9 
3 1 2 18 
7 1 2 3 20 9 18 9 
62 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
27 1 2 3 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 16 22 22 22 14 13 12 15 16 
27 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
15 1 2 3 4 6 5 7 8 9 10 10 10 10 17 19 
29 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 11 10 18 21 16 
3 1 2 18 
49 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 14 13 12 15 22 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
6 1 2 3 20 19 9 
17 1 2 3 9 4 6 5 7 8 9 11 10 13 14 15 12 16 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
16 1 2 3 20 4 6 5 7 8 9 11 10 16 18 21 16 
14 1 2 3 20 9 4 5 6 7 8 9 17 19 10 
3 1 2 18 
3 1 2 18 
17 1 2 3 9 9 9 4 5 6 7 8 9 10 10 17 19 10 
24 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
26 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
36 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
36 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 16 16 5 17 7 8 22 22 22 22 22 22 22 22 22 22 13 15 12 14 22 
30 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 15 13 12 14 16 
25 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 16 16 16 16 12 14 13 15 16 
29 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 12 14 13 15 16 
5 1 2 3 18 9 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
75 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 17 5 7 8 10 10 10 10 10 10 10 5 17 7 8 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 11 10 16 16 16 16 22 22 22 16 16 16 16 16 16 16 16 13 15 14 12 16 
3 1 2 18 
3 1 2 18 
34 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 21 18 16 
4 1 2 18 20 
4 1 2 18 20 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 14 12 15 13 16 
3 1 2 18 
25 1 2 3 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 14 13 12 15 22 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 13 14 15 12 16 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
22 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
38 1 2 3 9 4 5 6 7 8 9 10 10 17 5 7 8 10 11 10 16 22 22 22 5 17 7 8 22 22 22 11 22 16 14 12 15 13 16 
27 1 2 3 9 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 11 10 12 14 13 15 16 
7 1 2 3 4 9 18 9 
16 1 2 3 4 5 6 7 8 9 11 10 14 12 15 13 16 
3 1 2 18 
7 1 2 3 20 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
12 1 2 20 3 20 9 9 9 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
67 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 17 5 7 8 16 22 22 17 5 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 16 16 22 22 22 16 17 5 7 8 22 22 22 22 11 22 16 13 14 15 12 16 
4 1 2 18 20 
8 1 2 3 20 9 9 19 9 
22 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 11 10 15 13 12 14 16 
19 1 2 3 9 9 9 4 5 6 7 8 9 11 10 14 12 13 15 16 
21 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 9 9 19 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
22 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
3 1 2 18 
36 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
3 1 2 18 
23 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 16 16 22 17 19 22 
3 1 2 18 
3 1 2 18 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 17 19 10 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 19 9 
9 1 2 3 20 9 9 9 19 9 
9 1 2 20 20 3 20 9 18 9 
4 1 2 18 20 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 19 9 
29 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 16 22 22 22 22 13 12 14 15 16 
7 1 2 20 3 20 18 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
13 1 2 3 9 4 5 6 7 8 9 17 19 10 
4 1 2 18 20 
29 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 21 18 22 
6 1 2 3 20 18 9 
6 1 2 3 20 18 9 
4 1 2 18 20 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
25 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 16 16 16 22 22 15 13 14 12 16 
20 1 2 3 9 9 9 4 6 5 7 8 9 11 10 16 14 15 13 12 16 
6 1 2 3 20 18 9 
24 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 18 21 16 
41 1 2 20 3 20 9 4 5 6 7 8 9 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 13 14 15 12 16 
3 1 2 18 
38 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
12 1 2 3 4 6 5 7 8 9 19 17 10 
4 1 2 18 20 
21 1 2 3 4 5 6 7 8 9 11 10 16 16 16 22 22 12 14 15 13 16 
6 1 2 3 4 19 9 
22 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 17 19 10 
32 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
24 1 2 3 9 9 9 9 4 6 5 7 8 9 10 11 10 16 16 22 12 14 13 15 16 
22 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
27 1 2 3 9 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 16 14 13 15 12 16 
3 1 2 18 
6 1 2 3 20 18 9 
20 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 14 15 13 12 16 
39 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 16 16 22 22 17 5 7 8 22 22 22 11 22 16 14 15 13 12 22 
3 1 2 18 
29 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 12 14 15 13 16 
4 1 2 18 20 
23 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
40 1 2 3 9 4 6 5 7 8 9 10 10 10 10 11 10 17 5 7 8 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 18 21 16 
13 1 2 20 3 20 9 9 9 9 9 9 19 9 
4 1 2 18 20 
19 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
11 1 2 20 20 20 20 20 20 20 18 20 
16 1 2 3 9 9 4 6 5 7 8 9 10 10 19 17 10 
37 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 16 22 22 22 22 22 22 22 5 17 7 8 16 22 14 12 13 15 22 
17 1 2 3 4 5 6 7 8 9 11 10 16 14 13 12 15 16 
17 1 2 3 9 4 5 6 7 8 9 10 11 10 16 21 18 16 
3 1 2 18 
14 1 2 3 4 6 5 7 8 9 11 10 18 21 16 
47 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 16 16 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 21 18 16 
6 1 2 3 20 18 9 
23 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 21 18 16 
27 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
31 1 2 3 9 9 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 11 10 16 22 22 22 12 14 13 15 16 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 15 13 12 16 
32 1 2 3 20 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 18 21 16 
12 1 2 3 9 9 9 9 9 9 9 9 19 
23 1 2 3 20 4 6 5 7 8 9 10 11 10 16 16 22 22 22 14 13 12 15 16 
3 1 2 18 
17 1 2 3 9 4 6 5 7 8 9 11 10 15 12 14 13 16 
8 1 2 3 9 9 9 19 9 
36 1 2 3 20 4 9 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 5 17 7 8 10 10 11 10 16 16 22 22 21 18 22 
3 1 2 18 
5 1 2 20 18 20 
8 1 2 3 9 9 9 18 9 
21 1 2 3 4 5 6 7 8 9 11 10 16 16 16 22 22 13 14 15 12 16 
7 1 2 3 20 9 19 9 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
28 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 16 22 22 22 22 13 12 14 15 16 
3 1 2 18 
16 1 2 3 20 9 4 6 5 7 8 9 11 10 21 18 16 
4 1 2 18 20 
6 1 2 3 9 19 9 
30 1 2 3 20 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 16 22 22 13 14 15 12 22 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 9 
8 1 2 3 20 9 9 18 9 
17 1 2 3 9 4 6 5 7 8 9 11 10 14 13 12 15 16 
12 1 2 3 20 9 9 9 9 9 9 19 9 
23 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
5 1 2 3 19 9 
4 1 2 18 20 
31 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 11 10 14 15 12 13 16 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 14 12 13 15 16 
15 1 2 3 4 5 6 7 8 9 10 11 10 18 21 16 
43 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 11 10 16 14 13 12 15 16 
3 1 2 18 
42 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
23 1 2 3 9 9 9 9 4 6 5 7 8 9 10 11 10 16 16 16 16 18 21 16 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 12 14 13 15 16 
21 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 14 12 13 15 16 
24 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
29 1 2 20 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
32 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 16 18 21 16 
18 1 2 3 20 4 5 6 7 8 9 11 10 16 13 14 12 15 16 
17 1 2 3 20 4 5 6 7 8 9 10 10 10 10 17 19 10 
22 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
40 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 14 13 15 12 16 
3 1 2 18 
17 1 2 3 20 4 5 6 7 8 9 11 10 13 14 12 15 16 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 12 13 15 16 
5 1 2 3 18 9 
6 1 2 3 20 18 9 
24 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 12 13 15 14 16 
4 1 2 18 20 
5 1 2 20 18 20 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 16 14 13 15 12 16 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 14 12 15 13 16 
16 1 2 3 9 4 6 5 7 8 9 10 10 10 10 19 17 
3 1 2 18 
31 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
34 1 2 3 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 16 5 17 7 8 16 14 13 15 12 22 
21 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 14 13 12 15 16 
22 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 16 18 21 16 
31 1 2 3 20 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 11 10 16 22 22 16 16 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
31 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
3 1 2 18 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 14 13 12 15 16 
23 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
17 1 2 3 9 9 9 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
26 1 2 3 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 11 10 21 18 16 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
6 1 2 3 20 18 9 
9 1 2 3 9 9 9 9 19 9 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 23 14 12 15 13 16 
36 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 11 10 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
5 1 2 23 18 23 
22 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
24 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
5 1 2 20 18 20 
5 1 2 20 18 20 
26 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 13 14 12 15 16 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 14 15 13 12 16 
5 1 2 23 18 23 
28 1 2 3 4 6 5 7 8 9 5 17 7 8 10 11 10 16 16 22 22 22 22 16 14 12 15 13 16 
28 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 5 17 7 8 16 13 14 12 15 22 
33 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 5 17 7 8 16 14 13 12 15 22 
14 1 2 3 9 9 9 9 9 9 9 9 9 19 9 
5 1 2 20 18 20 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 14 12 15 13 16 
3 1 2 18 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 12 14 15 13 16 
4 1 2 18 20 
27 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 16 22 22 18 21 22 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 18 21 16 
3 1 2 18 
27 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
33 1 2 3 20 4 6 5 7 8 9 5 17 7 8 10 10 10 10 11 10 16 22 16 5 17 7 8 16 15 14 12 13 22 
30 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
6 1 2 3 9 18 9 
23 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 12 14 13 15 16 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
28 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 14 12 13 15 16 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 18 21 16 
36 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 16 22 22 16 16 22 22 22 16 13 14 15 12 16 
11 1 2 3 9 9 9 9 9 9 9 19 
10 1 2 3 20 9 9 9 9 18 9 
8 1 2 3 20 9 9 18 9 
25 1 2 3 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 11 10 15 13 12 14 16 
3 1 2 18 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
52 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 17 5 7 8 22 22 22 22 22 22 11 22 16 22 22 22 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 21 18 22 
17 1 2 3 9 4 6 5 7 8 9 11 10 13 15 14 12 16 
19 1 2 3 9 9 4 5 6 7 8 9 10 11 10 13 14 12 15 16 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
31 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
7 1 2 3 4 9 19 9 
6 1 2 3 9 19 9 
30 1 2 3 9 9 9 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 16 16 16 14 12 13 15 16 
3 1 2 18 
7 1 2 3 20 9 18 9 
20 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 16 21 18 16 
5 1 2 20 18 20 
19 1 2 3 9 9 4 6 5 7 8 9 10 11 10 13 15 14 12 16 
15 1 2 3 4 5 6 7 8 9 10 10 10 19 17 10 
21 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 11 10 21 18 16 
23 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 22 22 22 14 15 13 12 16 
23 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 22 16 12 13 14 15 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 12 15 14 16 
9 1 2 3 20 9 9 9 18 9 
28 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 22 22 22 22 13 15 14 12 16 
27 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 22 14 15 13 12 16 
6 1 2 3 20 18 9 
49 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 22 11 22 14 12 13 15 16 
16 1 2 3 20 9 9 4 5 6 7 8 9 10 19 17 10 
7 1 2 3 9 9 19 9 
16 1 2 3 4 5 6 7 8 9 11 10 14 13 12 15 16 
4 1 2 18 20 
25 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
27 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 16 22 12 14 13 15 16 
35 1 2 3 9 9 4 6 5 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 11 10 16 14 13 15 12 16 
27 1 2 20 3 20 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 16 16 12 13 15 14 16 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
6 1 2 3 9 18 9 
18 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 19 17 10 
3 1 2 18 
9 1 2 3 9 9 9 9 9 19 
4 1 2 18 20 
5 1 2 3 18 9 
7 1 2 23 23 23 18 23 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
31 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 11 10 16 22 22 22 22 22 22 22 22 22 17 19 22 
16 1 2 3 20 4 6 5 7 8 9 10 11 10 18 21 16 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
24 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 16 16 23 16 14 15 12 13 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
25 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
17 1 2 3 9 9 4 5 6 7 8 9 11 10 16 21 18 16 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 15 14 13 12 16 
4 1 2 18 20 
34 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 11 10 16 16 13 12 14 15 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
7 1 2 3 20 9 18 9 
38 1 2 3 9 9 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 16 22 22 22 22 21 18 16 
25 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 16 16 22 22 21 18 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
38 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 11 10 18 21 16 
39 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
22 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 22 16 14 12 13 15 16 
4 1 2 18 20 
23 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 13 14 15 12 16 
4 1 2 18 20 
6 1 2 3 20 18 9 
17 1 2 3 4 5 6 7 8 9 10 11 10 12 13 15 14 16 
4 1 2 18 20 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
14 1 2 3 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
29 1 2 3 4 6 5 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 14 15 13 12 16 
4 1 2 18 20 
18 1 2 3 9 9 4 5 6 7 8 9 11 10 13 14 12 15 16 
5 1 2 20 18 20 
4 1 2 18 20 
15 1 2 3 9 4 6 5 7 8 9 11 10 21 18 16 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
12 1 2 3 20 9 9 9 9 9 9 18 9 
30 1 2 20 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 11 10 14 13 12 15 16 
23 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 16 22 22 13 15 14 12 16 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 14 13 15 12 16 
6 1 2 3 20 18 9 
7 1 2 3 20 9 18 9 
29 1 2 3 4 6 5 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 12 13 15 14 16 
27 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
9 1 2 3 9 9 9 9 18 9 
4 1 2 18 20 
21 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 22 14 13 12 15 16 
7 1 2 3 4 9 19 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
38 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 17 19 
32 1 2 3 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
19 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
23 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 22 22 22 14 13 15 12 16 
14 1 2 3 9 4 5 6 7 8 9 10 19 17 10 
28 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 19 17 22 
4 1 2 18 20 
12 1 2 3 20 9 9 9 9 9 9 19 9 
19 1 2 20 20 3 20 9 9 4 6 5 7 8 9 10 10 17 19 10 
18 1 2 3 20 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
35 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 17 19 10 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
41 1 2 3 20 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 16 22 22 14 15 13 12 16 
4 1 2 18 20 
24 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 18 21 16 
3 1 2 18 
30 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 16 14 13 12 15 16 
3 1 2 18 
7 1 2 3 9 9 19 9 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 13 12 15 16 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 21 18 16 
3 1 2 18 
35 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 16 16 22 22 22 22 16 22 22 22 22 22 22 22 14 13 12 15 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
29 1 2 3 20 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 11 10 16 16 16 14 15 13 12 16 
3 1 2 18 
42 1 2 3 20 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 16 5 17 7 8 16 13 12 14 15 22 
22 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
26 1 2 20 3 20 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 13 14 12 15 16 
23 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
10 1 2 3 9 9 9 9 9 9 19 
24 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 11 10 16 22 15 13 12 14 16 
19 1 2 3 20 4 5 6 7 8 9 10 11 10 16 14 12 13 15 16 
3 1 2 18 
43 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 21 18 16 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 19 17 
5 1 2 20 18 20 
5 1 2 3 19 9 
23 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 22 22 16 22 22 18 21 16 
38 1 2 3 20 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 16 13 14 12 15 16 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 14 12 13 15 16 
20 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 10 
6 1 2 3 9 19 9 
29 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 16 22 22 22 22 22 14 13 15 12 16 
20 1 2 20 3 20 4 5 6 7 8 9 10 17 5 7 8 10 17 19 10 
4 1 2 18 20 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
20 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 14 13 15 12 16 
27 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 16 22 22 12 13 14 15 16 
12 1 2 3 4 6 5 7 8 9 19 17 10 
3 1 2 18 
19 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
4 1 2 18 20 
23 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 16 22 22 15 13 12 14 16 
24 1 2 3 20 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 19 17 22 
3 1 2 18 
15 1 2 3 20 9 4 5 6 7 8 9 10 17 19 10 
28 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 22 22 22 22 12 13 14 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
7 1 2 3 20 9 18 9 
9 1 2 3 9 9 9 9 19 9 
7 1 2 3 9 9 9 19 
3 1 2 18 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 14 15 12 13 16 
9 1 2 20 20 20 3 20 18 9 
24 1 2 3 9 4 6 5 7 8 9 10 10 5 17 7 8 10 11 10 14 13 12 15 16 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
27 1 2 3 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 11 10 14 15 13 12 16 
3 1 2 18 
7 1 2 3 20 9 19 9 
5 1 2 20 18 20 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 19 17 
13 1 2 3 9 4 6 5 7 8 9 17 19 10 
6 1 2 3 20 18 9 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
5 1 2 3 19 9 
3 1 2 18 
32 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 11 10 16 16 22 22 22 16 14 15 13 12 16 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 15 14 12 13 16 
25 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 16 12 15 13 14 16 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 18 21 16 
12 1 2 3 20 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 14 12 13 15 16 
4 1 2 18 20 
33 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
5 1 2 3 19 9 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 14 13 12 15 16 
31 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 17 5 7 8 10 10 11 10 16 22 15 13 12 14 16 
6 1 2 20 20 18 20 
21 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 19 10 
8 1 2 3 9 9 9 19 9 
28 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 21 18 22 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
20 1 2 3 4 6 5 7 8 9 10 11 10 16 16 16 13 14 15 12 16 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
22 1 2 20 20 20 20 20 3 20 4 6 5 7 8 9 11 10 15 13 14 12 16 
19 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
38 1 2 20 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 5 17 7 8 10 11 10 16 22 5 17 7 8 22 22 22 22 21 18 22 
4 1 2 18 20 
24 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 16 13 14 15 12 16 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 3 19 9 
22 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
14 1 2 3 20 9 4 6 5 7 8 9 19 17 10 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
13 1 2 3 20 9 9 9 9 9 9 9 19 9 
28 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 16 13 14 15 12 16 
15 1 2 3 20 9 4 6 5 7 8 9 10 17 19 10 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
4 1 2 18 20 
19 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 10 19 17 10 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
5 1 2 20 18 20 
3 1 2 18 
6 1 2 3 20 19 9 
10 1 2 3 20 9 9 9 9 18 9 
5 1 2 3 19 9 
22 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 17 19 10 
3 1 2 18 
24 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
46 1 2 3 9 4 5 6 7 8 9 10 10 11 10 17 5 7 8 16 22 22 22 22 5 17 7 8 22 22 22 22 22 22 11 22 16 5 17 7 8 16 14 12 13 15 22 
4 1 2 18 20 
26 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 14 12 13 15 16 
23 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
9 1 2 3 9 9 9 9 18 9 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 11 10 16 16 16 16 22 13 14 15 12 16 
11 1 2 3 20 9 9 9 9 9 19 9 
3 1 2 18 
8 1 2 20 20 3 20 19 9 
6 1 2 3 20 18 9 
6 1 2 3 9 18 9 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
3 1 2 18 
25 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
4 1 2 18 20 
14 1 2 3 9 9 4 6 5 7 8 9 10 19 17 
25 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 12 14 15 13 16 
25 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 11 10 14 13 12 15 16 
29 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
23 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 19 17 10 
4 1 2 18 20 
16 1 2 3 20 4 5 6 7 8 9 10 11 10 21 18 16 
3 1 2 18 
6 1 2 3 9 18 9 
22 1 2 3 4 6 5 7 8 9 10 11 10 16 16 22 22 22 14 13 12 15 16 
17 1 2 3 9 4 6 5 7 8 9 10 10 11 10 18 21 16 
3 1 2 18 
7 1 2 3 9 9 18 9 
19 1 2 3 9 9 4 5 6 7 8 9 10 11 10 13 14 15 12 16 
5 1 2 20 18 20 
14 1 2 20 3 20 9 9 9 9 9 9 9 18 9 
18 1 2 3 20 9 4 6 5 7 8 9 11 10 15 13 12 14 16 
4 1 2 18 20 
19 1 2 3 4 6 5 7 8 9 11 10 16 22 22 13 12 14 15 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 19 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 17 19 22 
4 1 2 18 20 
4 1 2 18 20 
40 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 22 16 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 11 22 14 13 12 15 16 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 9 4 5 6 7 8 9 10 11 10 16 21 18 16 
21 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 19 10 
16 1 2 3 4 5 6 7 8 9 10 11 10 16 17 19 16 
4 1 2 18 20 
3 1 2 18 
10 1 2 20 3 20 9 9 9 18 9 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
4 1 2 18 20 
13 1 2 3 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 19 9 
3 1 2 18 
6 1 2 3 9 18 9 
3 1 2 18 
13 1 2 3 4 6 5 7 8 9 10 18 21 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
19 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
19 1 2 3 4 6 5 7 8 9 10 11 10 16 16 13 14 12 15 16 
12 1 2 3 4 5 6 7 8 9 17 19 10 
6 1 2 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
5 1 2 20 18 20 
16 1 2 3 4 5 6 7 8 9 10 10 11 10 21 18 16 
32 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 23 23 16 22 22 22 22 22 22 22 22 22 16 18 21 16 
24 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 13 14 12 15 16 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 21 18 16 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
30 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
14 1 2 3 9 4 6 5 7 8 9 10 17 19 10 
5 1 2 3 18 9 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 12 13 15 14 16 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 19 17 10 
16 1 2 3 20 4 5 6 7 8 9 10 10 10 10 19 17 
3 1 2 18 
21 1 2 3 20 9 9 4 6 5 7 8 9 10 11 10 16 16 16 21 18 16 
3 1 2 18 
13 1 2 3 20 4 5 6 7 8 9 17 19 10 
22 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 14 15 13 12 16 
18 1 2 3 9 9 4 5 6 7 8 9 11 10 14 13 12 15 16 
4 1 2 18 20 
10 1 2 3 20 9 9 9 9 18 9 
16 1 2 3 9 4 6 5 7 8 9 10 10 10 17 19 10 
16 1 2 3 4 6 5 7 8 9 11 10 13 14 12 15 16 
7 1 2 3 20 9 18 9 
19 1 2 3 9 9 4 6 5 7 8 9 10 11 10 13 14 15 12 16 
20 1 2 3 4 5 6 7 8 9 11 10 16 16 16 16 13 15 12 14 16 
4 1 2 18 20 
11 1 2 3 20 4 9 9 9 9 19 9 
25 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
14 1 2 3 20 9 9 9 9 9 9 9 9 18 9 
28 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 13 14 12 15 16 
30 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 22 13 12 14 15 16 
34 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 11 10 16 16 22 22 22 22 22 13 14 15 12 16 
11 1 2 3 20 9 9 9 9 9 18 9 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
30 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
26 1 2 3 9 9 4 5 6 7 8 9 10 10 5 17 7 8 10 10 11 10 14 12 13 15 16 
11 1 2 3 9 9 9 9 9 9 19 9 
3 1 2 18 
14 1 2 3 20 9 4 5 6 7 8 9 17 19 10 
22 1 2 20 3 20 4 5 6 7 8 9 10 10 10 10 11 10 14 15 13 12 16 
37 1 2 3 4 6 5 7 8 9 11 10 16 16 16 22 22 22 22 22 22 16 16 16 16 16 16 16 16 16 22 22 22 13 14 15 12 16 
16 1 2 3 4 6 5 7 8 9 11 10 14 12 15 13 16 
4 1 2 18 20 
4 1 2 18 20 
34 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 10 17 
8 1 2 3 9 9 9 19 9 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 15 13 12 16 
4 1 2 18 20 
18 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
21 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 16 16 21 18 16 
7 1 2 3 9 9 19 9 
3 1 2 18 
32 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 14 13 15 12 16 
22 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
35 1 2 3 4 6 5 7 8 9 10 10 17 5 7 8 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 19 17 10 
15 1 2 3 9 4 6 5 7 8 9 11 10 18 21 16 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
6 1 2 3 9 18 9 
3 1 2 18 
3 1 2 18 
21 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 17 19 10 
11 1 2 3 9 9 9 9 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
45 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 14 12 13 15 16 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 10 10 11 10 21 18 16 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
6 1 2 3 9 18 9 
3 1 2 18 
5 1 2 20 18 20 
27 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 16 14 13 15 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 13 12 15 16 
25 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 21 18 16 
4 1 2 18 20 
40 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 16 14 15 13 12 16 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
27 1 2 3 4 5 6 7 8 9 5 17 7 8 10 17 5 7 8 10 10 10 10 10 10 10 19 17 
30 1 2 3 20 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 18 21 16 
33 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 16 22 19 17 22 
44 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 5 17 7 8 16 22 22 22 22 22 22 22 22 22 11 22 16 22 22 13 14 12 15 16 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 9 19 9 
11 1 2 3 20 9 9 9 9 9 18 9 
28 1 2 3 20 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 17 19 10 
10 1 2 20 20 3 20 9 9 18 9 
3 1 2 18 
10 1 2 3 20 9 9 9 9 19 9 
8 1 2 3 9 9 9 18 9 
9 1 2 20 20 3 20 9 19 9 
18 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 17 19 10 
32 1 2 23 23 20 23 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 22 14 12 13 15 16 
4 1 2 18 20 
22 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 9 
31 1 2 3 4 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 5 17 7 8 10 10 10 10 10 19 17 10 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
28 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 11 10 16 18 21 16 
17 1 2 3 20 9 9 9 4 5 6 7 8 9 10 19 17 10 
30 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 16 5 17 7 8 16 22 22 19 17 22 
3 1 2 18 
58 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 17 19 22 
27 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 22 22 16 16 15 13 14 12 16 
25 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 16 16 22 22 22 16 21 18 16 
19 1 2 3 4 6 5 7 8 9 10 11 10 16 22 15 13 14 12 16 
17 1 2 3 20 4 6 5 7 8 9 11 10 13 14 15 12 16 
18 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 21 18 16 
8 1 2 3 20 9 4 19 9 
3 1 2 18 
23 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 16 22 22 16 16 21 18 16 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 9 9 4 6 5 7 8 9 10 11 10 12 13 15 14 16 
4 1 2 18 20 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 21 18 16 
3 1 2 18 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 11 10 19 17 16 
5 1 2 3 19 9 
4 1 2 18 20 
20 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 14 13 12 15 16 
6 1 2 3 20 18 9 
3 1 2 18 
70 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 5 17 7 8 22 22 22 22 22 22 11 22 13 14 15 12 16 
4 1 2 18 20 
5 1 2 20 18 20 
3 1 2 18 
23 1 2 3 20 9 9 9 9 9 4 6 5 7 8 9 10 11 10 14 12 13 15 16 
8 1 2 3 9 9 9 18 9 
3 1 2 18 
27 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 16 16 16 16 16 22 22 14 13 12 15 16 
8 1 2 3 9 9 9 19 9 
4 1 2 18 20 
28 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
30 1 2 3 9 9 4 5 6 7 8 9 11 10 17 5 7 8 16 22 22 22 22 22 11 22 14 15 13 12 16 
20 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
19 1 2 3 20 9 9 9 9 4 5 6 7 8 9 11 10 18 21 16 
4 1 2 18 20 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
39 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 16 22 22 22 16 16 22 22 22 16 16 16 16 16 22 22 22 22 22 14 15 13 12 16 
3 1 2 18 
21 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 17 19 10 
5 1 2 20 18 20 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 9 9 9 
4 1 2 18 20 
35 1 2 3 20 9 4 9 9 9 9 9 9 9 9 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 11 10 21 18 16 
3 1 2 18 
40 1 2 3 20 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 11 10 16 22 22 17 19 22 
65 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 14 15 13 12 22 
25 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 13 15 12 14 16 
4 1 2 18 20 
5 1 2 3 18 9 
3 1 2 18 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
6 1 2 3 20 18 9 
45 1 2 3 20 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 16 13 14 12 15 16 
4 1 2 18 20 
12 1 2 3 9 9 9 9 9 9 9 19 9 
24 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 17 19 22 
8 1 2 20 3 20 9 18 9 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 14 15 13 12 16 
4 1 2 18 20 
3 1 2 18 
26 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 13 14 15 12 16 
24 1 2 3 9 9 4 6 5 7 8 9 11 10 16 22 22 22 22 16 14 12 13 15 16 
5 1 2 23 18 23 
6 1 2 3 20 18 9 
5 1 2 3 18 9 
24 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
37 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 19 17 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 13 14 12 15 16 
4 1 2 18 20 
6 1 2 3 20 18 9 
4 1 2 18 20 
6 1 2 20 20 18 20 
3 1 2 18 
19 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
3 1 2 18 
16 1 2 3 9 9 9 4 6 5 7 8 9 10 17 19 10 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 14 12 13 15 16 
6 1 2 3 9 18 9 
3 1 2 18 
26 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
10 1 2 3 20 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
27 1 2 3 9 9 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 11 10 14 15 13 12 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
28 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 22 22 16 22 22 22 22 22 14 13 15 12 16 
4 1 2 18 20 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 14 13 15 12 16 
3 1 2 18 
19 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
6 1 2 3 9 18 9 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 16 21 18 16 
24 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
45 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 18 21 22 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 13 14 15 12 16 
3 1 2 18 
5 1 2 20 18 20 
5 1 2 20 18 20 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
3 1 2 18 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
17 1 2 3 9 9 9 9 4 5 6 7 8 9 10 17 19 10 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 17 19 10 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 13 12 15 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
11 1 2 20 3 20 9 9 9 4 18 9 
25 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 19 17 10 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 17 19 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
9 1 2 3 9 9 9 9 9 19 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 12 13 15 16 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
15 1 2 3 9 4 5 6 7 8 9 10 10 19 17 10 
32 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 16 22 16 5 17 7 8 16 14 13 15 12 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 9 4 6 5 7 8 9 11 10 14 15 13 12 16 
22 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 14 12 15 13 16 
22 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 22 16 14 13 12 15 16 
44 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 5 17 7 8 10 10 10 10 10 10 11 10 16 5 17 7 8 16 22 22 22 22 22 14 15 13 12 22 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 16 18 21 16 
3 1 2 18 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
18 1 2 20 3 20 9 4 6 5 7 8 9 11 10 16 21 18 16 
22 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 10 17 
16 1 2 3 9 9 4 5 6 7 8 9 10 10 19 17 10 
20 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 13 14 12 15 16 
31 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 16 5 17 7 8 22 22 22 11 22 15 13 12 14 16 
4 1 2 18 20 
22 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 16 16 14 12 15 13 16 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
19 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
30 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 17 19 
22 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 11 10 13 14 12 15 16 
29 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 16 22 22 15 14 13 12 16 
3 1 2 18 
15 1 2 3 9 9 4 6 5 7 8 9 10 19 17 10 
4 1 2 18 20 
31 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 16 22 22 22 22 13 14 15 12 22 
14 1 2 3 20 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 11 10 13 12 14 15 16 
7 1 2 3 9 4 19 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
27 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 16 22 22 22 22 22 22 22 22 17 19 22 
4 1 2 18 20 
25 1 2 3 20 4 5 6 7 8 9 11 10 16 16 22 22 22 22 22 22 13 14 12 15 16 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 11 10 13 14 15 12 16 
4 1 2 18 20 
20 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
5 1 2 20 18 20 
6 1 2 3 20 19 9 
3 1 2 18 
3 1 2 18 
27 1 2 3 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 16 14 15 13 12 16 
23 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 14 12 15 13 16 
34 1 2 3 20 4 6 5 7 8 9 10 5 17 7 8 10 17 5 7 8 10 17 5 7 8 10 11 10 16 14 12 13 15 16 
26 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 22 13 15 12 14 16 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 17 19 10 
5 1 2 3 18 9 
4 1 2 18 20 
22 1 2 3 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 19 17 10 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 13 12 14 15 16 
31 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 16 22 22 12 13 15 14 16 
24 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
22 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 17 19 
3 1 2 18 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 10 
20 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 11 10 21 18 16 
11 1 2 3 20 9 9 9 9 9 18 9 
20 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 11 10 21 18 16 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 12 14 13 15 16 
3 1 2 18 
3 1 2 18 
24 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 14 13 15 12 16 
4 1 2 18 20 
16 1 2 3 4 6 5 7 8 9 11 10 14 12 13 15 16 
4 1 2 18 20 
6 1 2 3 20 18 9 
44 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 19 10 17 
3 1 2 18 
6 1 2 3 9 19 9 
4 1 2 18 20 
3 1 2 18 
41 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 11 22 14 15 13 12 16 
3 1 2 18 
8 1 2 3 9 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
20 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 21 18 16 
3 1 2 18 
3 1 2 18 
53 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 16 17 5 7 8 16 22 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 11 22 12 13 15 14 16 
3 1 2 18 
62 1 2 3 20 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 11 10 16 5 17 7 8 16 22 22 22 22 22 22 22 22 15 13 12 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 
7 1 2 3 9 4 19 9 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 14 15 12 16 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
6 1 2 3 20 18 9 
4 1 2 18 20 
17 1 2 3 20 4 5 6 7 8 9 10 10 11 10 21 18 16 
24 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
44 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 16 16 14 13 12 15 16 
8 1 2 3 9 9 4 19 9 
27 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 13 12 14 15 16 
6 1 2 3 20 18 9 
3 1 2 18 
36 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 14 13 12 15 16 
9 1 2 3 9 9 9 9 19 9 
11 1 2 3 20 9 9 9 9 9 18 9 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
14 1 2 3 20 9 9 9 9 9 9 9 9 19 9 
23 1 2 3 9 4 6 5 7 8 9 10 10 10 17 5 7 8 10 10 10 19 17 10 
20 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 13 14 12 15 16 
3 1 2 18 
6 1 2 3 9 19 9 
3 1 2 18 
8 1 2 3 9 9 4 18 9 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 17 19 10 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 12 13 15 16 
25 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 14 12 13 15 16 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 12 14 13 15 16 
21 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
5 1 2 3 19 9 
43 1 2 3 20 9 9 9 9 9 9 9 9 9 23 23 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 17 5 7 8 16 14 13 15 12 22 
20 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 13 14 12 15 16 
12 1 2 3 4 6 5 7 8 9 17 19 10 
14 1 2 3 20 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
33 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 10 11 10 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
16 1 2 3 9 9 4 5 6 7 8 9 10 10 17 19 10 
3 1 2 18 
5 1 2 3 19 9 
8 1 2 3 9 9 9 19 9 
19 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 19 17 10 
27 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 16 16 18 21 16 
3 1 2 18 
3 1 2 18 
33 1 2 3 20 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 5 17 7 8 16 13 15 14 12 22 
4 1 2 18 20 
14 1 2 3 20 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
26 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 14 12 13 15 16 
7 1 2 3 20 9 18 9 
3 1 2 18 
21 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 17 19 10 
3 1 2 18 
31 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 17 5 7 8 22 22 22 11 22 15 14 13 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 10 10 11 10 14 13 15 12 16 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 15 13 12 14 16 
33 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 17 5 7 8 10 11 10 16 22 16 16 22 22 13 14 15 12 16 
21 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 14 13 12 15 16 
27 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 14 13 15 12 16 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
16 1 2 3 9 9 4 5 6 7 8 9 10 10 17 19 10 
8 1 2 3 9 9 9 18 9 
3 1 2 18 
7 1 2 3 20 9 9 19 
3 1 2 18 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 22 14 12 13 15 16 
6 1 2 3 9 19 9 
8 1 2 3 9 9 9 9 19 
4 1 2 18 20 
22 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
27 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 13 14 15 12 16 
3 1 2 18 
4 1 2 18 20 
11 1 2 20 3 20 9 9 9 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 20 18 9 
25 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
21 1 2 3 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 19 17 10 
25 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 14 13 12 15 16 
3 1 2 18 
23 1 2 3 4 6 5 7 8 9 17 5 7 8 10 17 5 7 8 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
9 1 2 3 9 9 9 9 18 9 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
23 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 19 17 10 
17 1 2 3 9 9 4 6 5 7 8 9 10 11 10 18 21 16 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
47 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 5 17 7 8 10 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 14 13 15 12 16 
3 1 2 18 
31 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 16 22 22 22 17 19 22 
4 1 2 18 20 
3 1 2 18 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
19 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 18 21 16 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 18 9 
11 1 2 20 20 20 20 3 20 9 19 9 
10 1 2 20 3 20 9 9 9 18 9 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 19 17 10 
37 1 2 3 20 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 16 16 16 22 22 22 22 22 22 16 16 16 21 18 16 
3 1 2 18 
13 1 2 3 9 4 5 6 7 8 9 17 19 10 
4 1 2 18 20 
63 1 2 20 3 20 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 17 19 10 
32 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 17 5 7 8 22 22 22 11 22 12 13 15 14 16 
19 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 17 19 10 
27 1 2 3 9 4 5 6 7 8 9 11 10 16 16 16 22 22 22 22 22 16 16 14 13 12 15 16 
14 1 2 3 20 4 6 5 7 8 9 10 19 17 10 
21 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 21 18 16 
5 1 2 20 18 20 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
27 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
13 1 2 3 20 4 5 6 7 8 9 17 19 10 
19 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
8 1 2 3 20 9 9 18 9 
5 1 2 20 18 20 
25 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 14 12 13 15 16 
23 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 11 10 13 14 15 12 16 
3 1 2 18 
4 1 2 18 20 
10 1 2 20 20 3 20 9 9 18 9 
4 1 2 18 20 
30 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 16 16 22 22 22 16 14 15 13 12 16 
14 1 2 3 9 9 4 5 6 7 8 9 21 18 10 
18 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 18 21 16 
3 1 2 18 
5 1 2 3 18 9 
18 1 2 3 4 5 6 7 8 9 11 10 16 16 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
32 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 16 22 22 22 22 22 16 16 14 13 15 12 16 
31 1 2 3 4 5 6 7 8 9 10 11 10 16 5 17 7 8 22 17 5 7 8 22 22 11 22 14 12 13 15 16 
7 1 2 20 3 20 18 9 
21 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 16 13 14 15 12 16 
3 1 2 18 
3 1 2 18 
36 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 11 10 16 22 22 22 15 13 12 14 16 
4 1 2 18 20 
53 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 11 10 5 17 7 8 16 22 22 22 22 22 22 22 22 22 22 22 22 11 22 16 16 22 22 17 5 7 8 22 19 17 22 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 18 9 
22 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 16 14 15 13 12 16 
3 1 2 18 
3 1 2 18 
19 1 2 3 20 9 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
3 1 2 18 
28 1 2 3 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 13 15 12 16 
4 1 2 18 20 
26 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 14 12 13 15 16 
18 1 2 3 4 5 6 7 8 9 11 10 16 22 14 13 12 15 16 
28 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 11 10 16 16 16 14 12 13 15 16 
5 1 2 20 18 20 
40 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 16 5 17 7 8 22 22 22 22 22 22 22 22 11 22 13 14 15 12 16 
4 1 2 18 20 
6 1 2 3 9 19 9 
3 1 2 18 
34 1 2 3 20 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 14 13 15 12 16 
28 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 17 5 7 8 10 10 10 11 10 21 18 16 
3 1 2 18 
17 1 2 20 3 20 4 5 6 7 8 9 10 10 10 10 19 17 
5 1 2 23 18 23 
23 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 14 13 15 12 16 
3 1 2 18 
6 1 2 3 9 9 19 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
14 1 2 3 9 9 4 6 5 7 8 9 17 19 10 
4 1 2 18 20 
5 1 2 3 18 9 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 13 15 14 12 16 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
15 1 2 3 20 4 5 6 7 8 9 11 10 21 18 16 
4 1 2 18 20 
6 1 2 3 9 18 9 
27 1 2 3 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 21 18 16 
4 1 2 18 20 
24 1 2 3 20 4 6 5 7 8 9 10 10 10 17 5 7 8 10 10 11 10 18 21 16 
3 1 2 18 
32 1 2 3 20 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 10 11 10 16 22 22 22 14 15 13 12 22 
8 1 2 3 9 9 9 19 9 
18 1 2 3 4 5 6 7 8 9 11 10 16 22 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
30 1 2 3 20 9 4 6 5 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 10 10 11 10 18 21 16 
9 1 2 3 9 9 9 9 9 19 
20 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 14 12 13 15 16 
28 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 22 22 22 16 22 14 15 12 13 16 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
30 1 2 3 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 16 22 22 22 18 21 22 
3 1 2 18 
21 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 11 10 21 18 16 
28 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
27 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 14 13 15 12 16 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 13 15 12 16 
3 1 2 18 
25 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 13 14 15 12 16 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 14 12 13 15 16 
4 1 2 18 20 
4 1 2 18 20 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
29 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 18 21 16 
3 1 2 18 
4 1 2 18 20 
6 1 2 20 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 15 13 12 14 16 
4 1 2 18 20 
31 1 2 3 20 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 10 10 10 10 11 10 16 14 12 13 15 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
28 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 14 12 15 13 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 19 9 
45 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 22 22 22 22 22 22 22 16 22 22 22 16 16 22 22 22 22 22 16 22 22 14 15 13 12 16 
4 1 2 18 20 
5 1 2 3 18 9 
3 1 2 18 
24 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 14 13 15 12 16 
6 1 2 3 9 18 9 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 16 14 15 13 12 16 
33 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
37 1 2 3 20 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 17 5 7 8 10 10 10 10 10 11 10 12 14 15 13 16 
27 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 22 22 18 21 16 
3 1 2 18 
3 1 2 18 
33 1 2 3 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 17 5 7 8 10 10 10 10 10 17 19 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
12 1 2 3 9 9 9 9 9 9 9 18 9 
3 1 2 18 
42 1 2 3 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 11 10 16 16 22 22 22 22 22 22 22 22 22 17 5 7 8 16 13 14 15 12 22 
28 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
22 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 15 13 12 14 16 
4 1 2 18 20 
6 1 2 3 20 18 9 
12 1 2 3 9 9 9 9 9 9 9 9 19 
5 1 2 3 18 9 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 18 9 
5 1 2 3 19 9 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 20 4 5 6 7 8 9 10 10 10 17 19 10 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
5 1 2 3 18 9 
30 1 2 3 20 4 6 5 7 8 9 10 10 5 17 7 8 10 5 17 7 8 10 10 10 11 10 16 21 18 16 
3 1 2 18 
4 1 2 18 20 
31 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 17 5 7 8 10 10 10 10 11 10 14 12 15 13 16 
25 1 2 23 23 23 20 20 23 23 23 23 20 20 20 20 20 20 20 20 20 20 20 20 18 20 
3 1 2 18 
13 1 2 3 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
28 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
8 1 2 20 3 20 4 18 9 
5 1 2 3 18 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
29 1 2 20 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
7 1 2 3 9 9 19 9 
16 1 2 3 20 9 9 4 6 5 7 8 9 10 19 17 10 
4 1 2 18 20 
8 1 2 20 3 20 9 18 9 
23 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 14 13 15 12 16 
4 1 2 18 20 
4 1 2 18 20 
30 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 10 10 10 11 10 16 12 15 13 14 16 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 13 14 12 15 16 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
28 1 2 3 20 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 16 22 22 18 21 16 
4 1 2 18 20 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 10 10 11 10 18 21 16 
3 1 2 18 
25 1 2 20 3 20 4 5 6 7 8 9 10 17 5 7 8 10 10 11 10 12 14 13 15 16 
11 1 2 3 20 9 9 9 9 9 18 9 
4 1 2 18 20 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 20 3 20 4 6 5 7 8 9 10 11 10 16 15 14 12 13 16 
32 1 2 3 9 4 5 6 7 8 9 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 17 19 22 
5 1 2 20 18 20 
3 1 2 18 
25 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 16 12 14 13 15 16 
16 1 2 3 4 5 6 7 8 9 11 10 13 14 12 15 16 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
16 1 2 3 4 6 5 7 8 9 11 10 14 13 15 12 16 
13 1 2 3 20 4 6 5 7 8 9 17 19 10 
20 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 19 17 
8 1 2 3 9 9 9 19 9 
24 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
37 1 2 3 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 22 22 22 5 17 7 8 16 14 15 12 13 22 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 4 6 5 7 8 9 11 10 13 14 15 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
43 1 2 3 4 6 5 7 8 9 10 10 10 17 5 7 8 10 17 5 7 8 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 16 13 14 15 12 16 
4 1 2 18 20 
20 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 14 13 12 15 16 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 11 10 21 18 16 
24 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
6 1 2 3 9 19 9 
3 1 2 18 
4 1 2 18 20 
30 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
6 1 2 3 20 18 9 
50 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
10 1 2 3 20 9 9 9 9 9 19 
5 1 2 3 18 9 
4 1 2 18 20 
47 1 2 3 20 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 10 
5 1 2 20 18 20 
6 1 2 3 20 18 9 
10 1 2 3 9 9 9 9 9 19 9 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 19 17 10 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
3 1 2 18 
5 1 2 3 18 9 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 14 15 12 13 16 
16 1 2 3 20 9 9 4 5 6 7 8 9 10 17 19 10 
23 1 2 3 4 5 6 7 8 9 11 10 16 16 17 5 7 8 22 22 22 17 19 22 
17 1 2 3 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
12 1 2 3 4 6 5 7 8 9 21 18 10 
5 1 2 20 18 20 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 21 18 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
7 1 2 23 23 23 18 23 
3 1 2 18 
31 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 11 10 14 12 13 15 16 
11 1 2 3 20 9 9 9 9 4 19 9 
3 1 2 18 
5 1 2 20 18 20 
32 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
7 1 2 3 20 4 18 9 
6 1 2 3 20 18 9 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
14 1 2 3 4 6 5 7 8 9 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
36 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 16 23 23 23 16 22 22 22 22 22 22 22 22 22 22 16 13 14 15 12 16 
21 1 2 3 4 6 5 7 8 9 11 10 16 22 22 16 16 14 12 13 15 16 
20 1 2 3 9 4 5 6 7 8 9 11 10 16 16 16 13 15 14 12 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
20 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 14 13 15 12 16 
5 1 2 23 18 23 
26 1 2 20 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
15 1 2 3 4 6 5 7 8 9 11 10 16 21 18 16 
3 1 2 18 
23 1 2 3 4 5 6 7 8 9 11 10 16 22 22 16 22 22 22 15 14 12 13 16 
3 1 2 18 
4 1 2 18 20 
7 1 2 3 9 9 19 9 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 17 19 
25 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 22 13 14 12 15 16 
4 1 2 18 20 
26 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
32 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 11 10 16 22 22 22 18 21 22 
15 1 2 3 4 6 5 7 8 9 10 11 10 21 18 16 
21 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 12 13 15 14 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 5 17 7 8 10 11 10 14 15 12 13 16 
3 1 2 18 
8 1 2 3 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 11 10 14 13 12 15 16 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
33 1 2 3 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 16 13 12 15 14 16 
4 1 2 18 20 
5 1 2 3 19 9 
3 1 2 18 
35 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 22 11 22 12 14 13 15 16 
16 1 2 3 4 6 5 7 8 9 11 10 12 13 14 15 16 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 20 4 5 6 7 8 9 11 10 16 16 16 16 22 22 16 18 21 16 
3 1 2 18 
4 1 2 18 20 
32 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 14 15 12 13 16 
43 1 2 3 20 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 14 13 15 12 16 
3 1 2 18 
29 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
13 1 2 3 9 4 5 6 7 8 9 21 18 10 
21 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 14 13 15 12 16 
4 1 2 18 20 
13 1 2 3 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 17 19 10 
19 1 2 3 4 5 6 7 8 9 11 10 16 22 22 12 13 15 14 16 
3 1 2 18 
23 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 14 13 15 12 16 
24 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 14 13 15 12 16 
37 1 2 3 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 5 17 7 8 16 22 22 22 22 12 13 14 15 22 
26 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 16 16 16 16 14 15 13 12 16 
4 1 2 18 20 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 19 17 10 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 22 14 12 13 15 16 
4 1 2 18 20 
14 1 2 3 20 9 4 5 6 7 8 9 17 19 10 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
40 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 16 15 14 12 13 16 
26 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 11 10 12 13 14 15 16 
29 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 17 5 7 8 22 22 11 22 14 13 15 12 16 
26 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 16 16 16 22 22 22 14 12 15 13 16 
4 1 2 18 20 
20 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 11 10 18 21 16 
4 1 2 18 20 
3 1 2 18 
16 1 2 3 20 4 5 6 7 8 9 10 11 10 21 18 16 
4 1 2 18 20 
34 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 11 10 17 5 7 8 16 13 12 14 15 22 
25 1 2 3 4 6 5 7 8 9 17 5 7 8 10 11 10 16 22 22 22 14 13 15 12 16 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
34 1 2 3 20 4 5 6 7 8 9 10 17 5 7 8 10 10 11 10 16 22 22 22 22 22 22 22 16 16 15 13 12 14 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
12 1 2 3 4 6 5 7 8 9 17 19 10 
4 1 2 18 20 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
36 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 22 22 22 17 5 7 8 22 22 22 22 11 22 14 13 15 12 16 
24 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 19 17 10 
42 1 2 3 20 4 5 6 7 8 9 10 5 17 7 8 10 5 17 7 8 10 11 10 17 5 7 8 16 22 22 22 22 22 22 22 11 22 14 12 13 15 16 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 16 22 22 12 14 13 15 16 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
41 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 11 22 16 13 14 12 15 16 
4 1 2 18 20 
23 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 16 14 13 12 15 16 
7 1 2 3 20 9 18 9 
5 1 2 20 18 20 
38 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
26 1 2 3 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 17 19 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
16 1 2 3 4 5 6 7 8 9 11 10 14 12 15 13 16 
4 1 2 18 20 
5 1 2 3 18 9 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 13 15 12 16 
19 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 17 19 10 
3 1 2 18 
17 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 18 9 
25 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 14 15 13 12 16 
24 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 16 16 22 22 22 18 21 16 
17 1 2 3 4 5 6 7 8 9 5 17 7 8 10 19 17 10 
19 1 2 20 3 20 9 9 9 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
39 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 16 16 16 22 22 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 14 12 13 15 16 
7 1 2 3 9 9 19 9 
16 1 2 3 20 9 4 5 6 7 8 9 10 10 17 19 10 
8 1 2 3 9 9 9 18 9 
40 1 2 3 9 4 6 5 7 8 9 11 10 16 16 22 22 22 22 22 22 16 22 16 22 22 22 22 22 22 22 22 22 22 22 22 14 15 13 12 16 
5 1 2 20 18 20 
6 1 2 20 20 18 20 
3 1 2 18 
26 1 2 3 9 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 13 14 15 12 16 
11 1 2 3 9 9 9 9 9 4 19 9 
3 1 2 18 
6 1 2 3 9 19 9 
17 1 2 3 9 4 6 5 7 8 9 11 10 14 13 12 15 16 
30 1 2 20 3 20 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
18 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
4 1 2 18 20 
9 1 2 3 20 9 9 9 18 9 
9 1 2 3 9 9 9 9 18 9 
23 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 14 13 15 12 16 
3 1 2 18 
6 1 2 3 20 19 9 
3 1 2 18 
9 1 2 3 20 9 9 9 9 19 
40 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 14 12 13 15 16 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 14 12 15 13 16 
3 1 2 18 
33 1 2 3 4 5 6 7 8 9 17 5 7 8 10 5 17 7 8 10 11 10 16 22 22 22 22 16 22 22 22 19 17 22 
30 1 2 3 9 4 6 5 7 8 9 10 10 5 17 7 8 10 10 5 17 7 8 10 11 10 12 14 15 13 16 
3 1 2 18 
5 1 2 3 18 9 
5 1 2 3 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
32 1 2 3 9 4 6 5 7 8 9 10 10 5 17 7 8 10 10 10 10 10 10 10 11 10 16 16 14 15 12 13 16 
12 1 2 3 4 5 6 7 8 9 17 19 10 
16 1 2 3 4 6 5 7 8 9 10 11 10 16 18 21 16 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
21 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 14 15 13 12 16 
5 1 2 3 19 9 
7 1 2 3 9 9 9 19 
20 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 21 18 16 
22 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 11 10 12 13 14 15 16 
6 1 2 3 9 19 9 
5 1 2 20 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 11 10 14 15 13 12 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
5 1 2 3 19 9 
27 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
8 1 2 3 9 9 9 18 9 
66 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 21 18 16 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 19 17 10 
20 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 14 13 15 12 16 
10 1 2 20 3 20 9 9 9 18 9 
3 1 2 18 
18 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 21 18 16 
21 1 2 3 20 9 4 6 5 7 8 9 11 10 16 22 22 14 12 13 15 16 
24 1 2 3 9 4 9 9 6 5 7 8 9 10 11 10 16 16 22 22 12 14 15 13 16 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 3 19 9 
4 1 2 18 20 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 13 14 15 12 16 
7 1 2 3 20 9 18 9 
3 1 2 18 
26 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 13 14 12 15 16 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 13 14 15 12 16 
6 1 2 20 20 18 20 
20 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 13 14 12 15 16 
27 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
21 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
7 1 2 3 9 9 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
15 1 2 3 20 9 9 4 6 5 7 8 9 19 17 10 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 19 17 10 
11 1 2 3 20 9 9 9 9 4 19 9 
18 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 11 10 13 15 14 12 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
35 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 14 13 12 15 16 
3 1 2 18 
18 1 2 3 9 9 9 9 4 5 6 7 8 9 11 10 17 19 16 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
40 1 2 3 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 5 17 7 8 10 10 11 10 16 17 5 7 8 16 13 14 12 15 22 
4 1 2 18 20 
18 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 19 17 10 
17 1 2 3 9 4 5 6 7 8 9 11 10 15 14 12 13 16 
29 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 11 10 14 12 13 15 16 
3 1 2 18 
25 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 16 16 13 14 12 15 16 
6 1 2 3 9 19 9 
9 1 2 3 9 9 9 9 19 9 
3 1 2 18 
18 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 18 21 16 
20 1 2 3 9 4 6 5 7 8 9 11 10 16 22 16 14 15 13 12 16 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 9 4 6 5 7 8 9 11 10 13 12 14 15 16 
24 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 14 12 15 13 16 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 15 13 12 16 
33 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 5 17 7 8 16 22 22 22 22 22 22 11 22 14 13 15 12 16 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 19 17 
3 1 2 18 
5 1 2 3 18 9 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 12 13 15 16 
25 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 13 15 12 14 16 
17 1 2 3 4 6 5 7 8 9 10 10 11 10 16 21 18 16 
7 1 2 3 20 9 18 9 
48 1 2 3 20 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 11 10 16 16 16 16 16 22 22 22 22 12 13 15 14 22 
64 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 16 22 22 22 16 16 22 22 5 17 7 8 22 17 5 7 8 22 22 22 22 11 22 16 22 22 22 22 22 22 22 22 22 22 22 22 15 12 14 13 16 
8 1 2 20 3 20 9 18 9 
25 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 17 19 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
46 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 16 22 22 16 16 16 16 16 16 22 16 16 16 16 16 16 16 16 16 16 16 16 14 13 12 15 16 
4 1 2 18 20 
23 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
25 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 10 10 10 21 18 10 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 19 9 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
9 1 2 3 9 9 9 9 19 9 
36 1 2 3 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 16 22 22 17 5 7 8 16 14 12 13 15 22 
28 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
17 1 2 3 9 4 6 5 7 8 9 11 10 14 13 15 12 16 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 9 4 5 6 7 8 9 11 10 16 12 13 14 15 16 
33 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 11 10 16 16 16 22 14 12 13 15 16 
7 1 2 3 20 9 18 9 
22 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 11 10 14 12 13 15 16 
6 1 2 3 9 18 9 
22 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 17 19 10 
24 1 2 3 9 4 5 6 7 8 9 10 10 17 5 7 8 10 11 10 14 13 15 12 16 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 18 9 
30 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 22 22 16 16 14 12 13 15 16 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 17 19 10 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
22 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 19 17 
6 1 2 3 9 19 9 
44 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 16 22 22 22 16 15 13 14 12 16 
4 1 2 18 20 
5 1 2 3 19 9 
3 1 2 18 
16 1 2 3 9 4 6 5 7 8 9 11 10 16 17 19 22 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 14 13 15 12 16 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
36 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 10 11 10 16 16 22 22 22 22 22 17 5 7 8 16 15 13 12 14 22 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 3 19 9 
30 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 15 13 12 14 16 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 14 13 12 15 16 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
18 1 2 3 4 6 5 7 8 9 11 10 16 22 14 13 12 15 16 
24 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
23 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 14 15 12 13 16 
9 1 2 3 20 9 9 9 18 9 
6 1 2 3 4 19 9 
15 1 2 3 9 9 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
20 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 14 15 13 12 16 
5 1 2 3 19 9 
33 1 2 3 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 11 10 5 17 7 8 16 14 13 15 12 22 
3 1 2 18 
55 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
53 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 17 19 
19 1 2 3 20 9 4 6 5 7 8 9 10 11 10 14 13 15 12 16 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 18 9 
24 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 17 5 7 8 10 10 19 17 10 
26 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
6 1 2 3 20 18 9 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 11 10 16 16 14 13 15 12 16 
6 1 2 3 9 19 9 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 15 12 13 16 
30 1 2 3 4 6 5 7 8 9 5 17 7 8 10 11 10 16 22 22 22 5 17 7 8 16 12 13 15 14 22 
5 1 2 20 18 20 
34 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 17 5 7 8 22 22 22 22 22 22 22 22 11 22 14 13 15 12 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
13 1 2 3 20 4 5 6 7 8 9 17 19 10 
11 1 2 20 3 20 9 9 9 9 9 19 
21 1 2 3 20 9 4 6 5 7 8 9 10 10 11 10 16 23 16 21 18 22 
20 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
13 1 2 20 3 20 9 9 9 9 9 9 19 9 
27 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 14 12 15 13 16 
31 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 13 14 15 12 16 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
13 1 2 3 9 9 9 9 9 9 9 9 18 9 
15 1 2 3 9 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
33 1 2 3 4 6 5 7 8 9 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
7 1 2 3 20 9 19 9 
3 1 2 18 
15 1 2 3 20 4 6 5 7 8 9 11 10 18 21 16 
15 1 2 3 4 6 5 7 8 9 11 10 16 18 21 16 
6 1 2 3 9 19 9 
22 1 2 3 4 6 5 7 8 9 10 10 10 5 17 7 8 10 10 10 17 19 10 
25 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 15 13 12 14 16 
3 1 2 18 
29 1 2 3 4 5 6 7 8 9 10 10 10 10 17 5 7 8 10 10 10 10 10 11 10 13 14 15 12 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
4 1 2 18 20 
3 1 2 18 
33 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
20 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
24 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 14 12 15 13 16 
8 1 2 3 20 9 4 19 9 
16 1 2 3 4 6 5 7 8 9 11 10 14 12 15 13 16 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 9 4 5 6 7 8 9 11 10 16 18 21 16 
3 1 2 18 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 18 9 
27 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 11 10 16 16 22 14 12 15 13 16 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 18 9 
19 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 17 19 10 
25 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 14 15 12 13 16 
3 1 2 18 
21 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 14 13 12 15 16 
5 1 2 20 18 20 
31 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 16 22 22 16 16 14 13 15 12 16 
10 1 2 20 3 20 9 9 9 18 9 
23 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 13 14 12 15 16 
39 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 16 22 16 13 12 14 15 16 
3 1 2 18 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 11 10 15 12 14 13 16 
3 1 2 18 
26 1 2 3 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
33 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 16 22 22 22 22 16 22 22 22 14 12 13 15 16 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 13 12 15 16 
24 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 14 12 13 15 16 
4 1 2 18 20 
3 1 2 18 
35 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 11 10 16 16 22 22 22 14 12 15 13 16 
9 1 2 3 9 9 9 9 9 19 
5 1 2 3 18 9 
53 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 11 10 17 5 7 8 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 16 16 14 13 15 12 16 
9 1 2 3 20 9 9 9 18 9 
31 1 2 3 20 4 6 5 7 8 9 11 10 16 23 5 17 7 8 16 22 22 22 22 11 22 16 14 12 15 13 16 
26 1 2 3 20 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 15 13 14 12 16 
5 1 2 3 18 9 
16 1 2 3 9 4 5 6 7 8 9 11 10 16 18 21 16 
3 1 2 18 
17 1 2 3 20 9 4 5 6 7 8 9 10 11 10 21 18 16 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
3 1 2 18 
6 1 2 3 20 18 9 
7 1 2 3 20 9 19 9 
26 1 2 20 3 20 4 5 6 7 8 9 10 5 17 7 8 10 10 11 10 16 14 15 13 12 16 
25 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 13 14 12 15 16 
19 1 2 3 4 5 6 7 8 9 10 10 11 10 16 14 13 12 15 16 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
18 1 2 3 9 9 9 9 4 6 5 7 8 9 11 10 21 18 16 
5 1 2 20 18 20 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 11 10 16 16 18 21 16 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 16 14 15 13 12 16 
4 1 2 18 20 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
5 1 2 20 18 20 
10 1 2 20 3 20 9 9 9 18 9 
10 1 2 3 9 9 9 9 9 19 9 
4 1 2 18 20 
7 1 2 3 9 9 18 9 
24 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 13 14 15 12 16 
23 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 11 10 16 18 21 16 
7 1 2 3 9 9 18 9 
4 1 2 18 20 
21 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 15 14 13 12 16 
3 1 2 18 
42 1 2 3 4 6 5 7 8 9 10 10 17 5 7 8 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 17 19 22 
4 1 2 18 20 
8 1 2 3 9 9 9 18 9 
29 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 5 17 7 8 22 22 22 11 22 13 14 15 12 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
29 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 16 22 22 22 22 22 14 12 15 13 16 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
25 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
28 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 11 10 16 13 15 14 12 16 
18 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 17 19 10 
12 1 2 3 20 9 9 9 9 9 9 9 19 
20 1 2 3 20 9 9 9 9 9 4 6 5 7 8 9 10 10 19 17 10 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
16 1 2 3 4 5 6 7 8 9 11 10 14 13 12 15 16 
37 1 2 3 9 4 6 5 7 8 9 11 10 16 16 22 22 22 5 17 7 8 22 5 17 7 8 22 22 22 22 11 22 16 16 18 21 16 
39 1 2 20 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 22 22 22 22 22 16 16 17 5 7 8 22 19 17 22 
3 1 2 18 
4 1 2 18 20 
24 1 2 3 9 4 6 5 7 8 9 10 10 17 5 7 8 10 11 10 13 15 14 12 16 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 18 21 16 
3 1 2 18 
4 1 2 18 20 
44 1 2 3 20 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 16 16 22 12 14 15 13 16 
26 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 18 21 16 
7 1 2 3 9 9 18 9 
6 1 2 3 20 18 9 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
24 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
7 1 2 3 9 9 18 9 
22 1 2 3 20 9 9 9 4 5 6 7 8 9 10 11 10 16 12 13 15 14 16 
7 1 2 23 23 23 18 23 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
37 1 2 3 9 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 17 19 10 
6 1 2 3 20 18 9 
20 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 14 12 15 13 16 
3 1 2 18 
7 1 2 3 20 9 18 9 
40 1 2 3 20 4 6 5 7 8 9 10 10 5 17 7 8 10 10 10 10 10 10 10 17 5 7 8 10 5 17 7 8 10 11 10 13 14 15 12 16 
11 1 2 23 23 23 23 23 23 23 18 23 
22 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 15 14 13 12 16 
3 1 2 18 
21 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
4 1 2 18 20 
33 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 16 22 22 22 22 22 22 14 13 15 12 16 
25 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 22 16 22 22 16 14 13 15 12 16 
3 1 2 18 
17 1 2 3 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
5 1 2 3 18 9 
21 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 16 13 15 12 14 16 
4 1 2 18 20 
5 1 2 20 18 20 
23 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 11 10 16 22 17 19 16 
16 1 2 3 4 5 6 7 8 9 11 10 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
22 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 17 19 10 
3 1 2 18 
8 1 2 20 20 3 20 18 9 
3 1 2 18 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
6 1 2 3 20 18 9 
4 1 2 18 20 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
19 1 2 3 20 4 6 5 7 8 9 10 11 10 16 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
28 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 17 5 7 8 10 10 11 10 16 16 18 21 16 
3 1 2 18 
25 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 14 15 13 12 16 
3 1 2 18 
29 1 2 3 4 6 5 7 8 9 10 11 10 16 16 22 22 22 16 22 22 22 22 22 22 13 14 15 12 16 
20 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 15 12 13 14 16 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
23 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 11 10 16 16 16 13 15 12 
26 1 2 3 4 6 5 7 8 9 11 10 16 23 16 22 22 22 22 22 22 22 14 15 12 13 16 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 11 10 16 16 22 22 22 13 14 12 15 16 
27 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 16 16 22 22 22 16 14 12 13 15 16 
5 1 2 20 18 20 
26 1 2 3 4 6 5 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 14 12 15 13 16 
17 1 2 3 20 4 6 5 7 8 9 11 10 14 13 12 15 16 
23 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 14 15 13 12 16 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 9 9 9 19 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 13 14 12 15 16 
31 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 22 22 16 16 22 22 22 13 14 15 12 16 
4 1 2 18 20 
3 1 2 18 
32 1 2 3 9 9 9 4 6 5 7 8 9 11 10 17 5 7 8 16 22 22 22 22 22 22 11 22 12 13 15 14 16 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 9 9 19 9 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 12 15 13 16 
16 1 2 3 4 5 6 7 8 9 10 11 10 16 21 18 16 
40 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 17 19 10 
14 1 2 3 9 9 4 5 6 7 8 9 21 18 10 
26 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 14 15 12 13 16 
25 1 2 3 20 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 12 13 15 14 16 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 18 9 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 12 13 15 14 16 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 9 19 
8 1 2 3 20 9 9 18 9 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
23 1 2 20 3 20 4 6 5 7 8 9 10 10 11 10 16 22 22 14 13 12 15 16 
25 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 18 21 16 
6 1 2 3 9 18 9 
20 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 12 14 13 15 16 
4 1 2 18 20 
23 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 22 16 16 14 12 13 15 16 
6 1 2 3 20 18 9 
24 1 2 3 20 9 9 9 9 9 9 9 9 4 5 6 7 8 9 11 10 16 18 21 16 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 19 17 10 
34 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 16 22 17 5 7 8 16 22 22 22 11 22 16 16 14 13 15 12 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 14 12 13 15 16 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 11 10 18 21 16 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
28 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 22 22 17 19 
8 1 2 20 3 20 9 18 9 
13 1 2 20 3 20 9 9 9 9 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
16 1 2 3 20 4 6 5 7 8 9 10 11 10 21 18 16 
6 1 2 3 20 18 9 
4 1 2 18 20 
4 1 2 18 20 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
22 1 2 3 9 4 6 5 7 8 9 10 5 17 7 8 10 10 11 10 18 21 16 
20 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 10 17 19 10 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
30 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 5 17 7 8 10 10 10 11 10 14 13 15 12 16 
53 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 5 17 7 8 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
26 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 18 21 16 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
17 1 2 3 20 4 5 6 7 8 9 11 10 14 15 12 13 16 
4 1 2 18 20 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
8 1 2 3 9 9 9 9 19 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
6 1 2 3 9 18 9 
18 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 21 18 10 
3 1 2 18 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 14 13 12 15 16 
27 1 2 3 20 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 22 14 13 12 15 16 
7 1 2 3 20 4 19 9 
14 1 2 3 4 5 6 7 8 9 11 10 18 21 16 
17 1 2 3 4 5 6 7 8 9 10 10 10 11 10 21 18 16 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 
3 1 2 18 
17 1 2 3 9 9 4 5 6 7 8 9 10 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 17 19 10 
3 1 2 18 
25 1 2 3 9 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 11 10 18 21 16 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 22 14 13 15 12 16 
3 1 2 18 
10 1 2 3 20 9 9 9 9 18 9 
23 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 11 10 13 14 12 15 16 
20 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 19 17 10 
39 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 19 17 22 
3 1 2 18 
6 1 2 3 20 19 9 
25 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 16 22 22 22 22 22 17 19 22 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
5 1 2 3 19 9 
3 1 2 18 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 14 12 15 13 16 
4 1 2 18 20 
23 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 18 21 16 
4 1 2 18 20 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 11 10 16 16 15 13 12 14 16 
3 1 2 18 
34 1 2 3 4 5 6 7 8 9 10 10 11 10 16 17 5 7 8 16 22 22 22 22 11 22 16 16 22 22 14 12 13 15 16 
24 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
28 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 16 22 22 22 19 17 22 
8 1 2 20 3 20 9 18 9 
17 1 2 3 9 9 9 4 6 5 7 8 9 10 10 17 19 10 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 16 21 18 16 
3 1 2 18 
3 1 2 18 
22 1 2 3 9 9 9 9 9 4 6 5 7 8 9 11 10 16 14 15 13 12 16 
5 1 2 20 18 20 
3 1 2 18 
15 1 2 3 9 9 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
31 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 17 5 7 8 16 14 13 15 12 22 
14 1 2 20 3 20 4 6 5 7 8 9 10 19 17 
18 1 2 3 9 9 4 5 6 7 8 9 11 10 14 13 12 15 16 
3 1 2 18 
6 1 2 3 20 18 9 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
21 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 11 10 18 21 16 
21 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 14 12 13 15 16 
3 1 2 18 
30 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
4 1 2 18 20 
27 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 16 16 16 18 21 16 
4 1 2 18 20 
38 1 2 3 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 16 16 16 22 22 22 22 14 12 13 15 16 
8 1 2 3 20 9 9 9 19 
3 1 2 18 
28 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 16 22 16 16 16 16 12 13 15 14 16 
41 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 16 16 5 17 7 8 22 22 22 22 11 22 16 22 16 16 14 15 13 12 16 
18 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 19 17 10 
4 1 2 18 20 
23 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
21 1 2 3 20 9 4 5 6 7 8 9 11 10 16 22 22 13 15 14 12 16 
3 1 2 18 
22 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
7 1 2 3 9 9 19 9 
7 1 2 3 9 9 19 9 
28 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
4 1 2 18 20 
3 1 2 18 
30 1 2 3 20 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 16 16 18 21 16 
3 1 2 18 
3 1 2 18 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 10 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
13 1 2 3 9 4 6 5 7 8 9 10 19 17 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
24 1 2 3 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 19 17 10 
5 1 2 3 18 9 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 17 5 7 8 10 19 17 10 
26 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 22 14 13 12 15 16 
12 1 2 3 4 6 5 7 8 9 19 17 10 
15 1 2 3 4 6 5 7 8 9 10 11 10 21 18 16 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 18 21 16 
3 1 2 18 
43 1 2 3 20 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
36 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 16 16 16 16 14 12 13 15 16 
7 1 2 20 3 20 18 9 
27 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 17 5 7 8 10 10 19 17 10 
5 1 2 3 18 9 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
25 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 11 10 16 16 16 12 14 15 13 22 
17 1 2 3 20 4 5 6 7 8 9 11 10 14 15 13 12 16 
3 1 2 18 
5 1 2 20 18 20 
29 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 16 21 18 16 
19 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 17 19 10 
7 1 2 3 20 9 18 9 
6 1 2 3 20 19 9 
8 1 2 3 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
32 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
21 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 13 14 12 15 16 
7 1 2 3 20 9 18 9 
3 1 2 18 
17 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 17 19 
3 1 2 18 
5 1 2 3 19 9 
10 1 2 3 9 9 9 9 9 19 9 
18 1 2 3 4 5 6 7 8 9 11 10 16 22 14 13 12 15 16 
23 1 2 20 3 20 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 17 19 
15 1 2 3 4 5 6 7 8 9 10 11 10 21 18 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
23 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 19 17 
33 1 2 3 4 5 6 7 8 9 5 17 7 8 10 5 17 7 8 10 10 5 17 7 8 10 10 10 10 10 10 10 19 17 
12 1 2 3 4 6 5 7 8 9 19 17 10 
14 1 2 3 4 6 5 7 8 9 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
17 1 2 20 3 20 4 5 6 7 8 9 10 10 10 17 19 10 
22 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 17 19 
4 1 2 18 20 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
5 1 2 3 18 9 
5 1 2 3 18 9 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
5 1 2 3 18 9 
4 1 2 18 20 
4 1 2 18 20 
46 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 11 22 16 14 12 13 15 16 
37 1 2 3 4 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 5 17 7 8 10 11 10 16 5 17 7 8 16 14 12 15 13 22 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 20 9 9 9 4 6 5 7 8 9 10 11 10 14 13 12 15 16 
3 1 2 18 
40 1 2 3 4 5 6 7 8 9 5 17 7 8 10 5 17 7 8 10 17 5 7 8 10 10 10 10 10 11 10 17 5 7 8 16 13 12 14 15 22 
19 1 2 3 9 4 5 6 7 8 9 10 11 10 16 12 15 13 14 16 
23 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 13 15 14 12 16 
4 1 2 18 20 
6 1 2 3 9 19 9 
4 1 2 18 20 
17 1 2 3 4 5 6 7 8 9 11 10 16 14 13 15 12 16 
10 1 2 3 9 9 9 9 9 19 9 
4 1 2 18 20 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
6 1 2 3 20 19 9 
3 1 2 18 
7 1 2 3 9 9 18 9 
22 1 2 3 20 9 4 5 6 7 8 9 11 10 16 22 22 16 14 12 13 15 16 
3 1 2 18 
22 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 21 18 22 
9 1 2 3 9 9 9 9 18 9 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 10 19 17 
10 1 2 3 20 9 9 9 9 19 9 
16 1 2 3 9 9 4 5 6 7 8 9 10 10 17 19 10 
3 1 2 18 
26 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 19 17 
16 1 2 3 4 6 5 7 8 9 11 10 14 13 12 15 16 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
16 1 2 3 20 4 5 6 7 8 9 10 11 10 21 18 16 
20 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 19 17 
16 1 2 20 3 20 4 6 5 7 8 9 10 10 19 17 10 
4 1 2 18 20 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
35 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 22 14 13 12 15 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
22 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
6 1 2 3 20 18 9 
23 1 2 3 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 17 19 10 
6 1 2 3 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
6 1 2 3 20 18 9 
25 1 2 3 20 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 18 21 16 
24 1 2 3 20 4 5 6 7 8 9 10 10 17 5 7 8 10 11 10 13 15 12 14 16 
4 1 2 18 20 
17 1 2 3 4 5 6 7 8 9 10 11 10 13 14 12 15 16 
3 1 2 18 
47 1 2 3 20 9 4 6 5 7 8 9 10 11 10 16 22 22 22 16 16 22 22 22 22 22 22 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 13 14 12 15 16 
20 1 2 3 9 4 5 6 7 8 9 11 10 16 16 22 22 22 22 19 17 
18 1 2 3 4 6 5 7 8 9 11 10 16 16 15 14 12 13 16 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
22 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 13 14 12 15 16 
7 1 2 3 9 9 18 9 
38 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 16 22 22 16 16 16 16 14 13 12 15 16 
8 1 2 3 9 9 9 19 9 
3 1 2 18 
5 1 2 20 18 20 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 14 13 15 12 16 
26 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
21 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 13 14 12 15 16 
6 1 2 3 20 18 9 
8 1 2 20 20 3 20 18 9 
28 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 16 15 14 12 13 16 
4 1 2 18 20 
29 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 22 16 21 18 16 
26 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 12 13 15 14 16 
4 1 2 18 20 
4 1 2 18 20 
23 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 13 14 15 12 16 
6 1 2 20 20 18 20 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 10 17 19 
4 1 2 18 20 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 19 17 10 
5 1 2 20 18 20 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 19 17 22 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
11 1 2 20 3 20 9 9 9 9 18 9 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
4 1 2 18 20 
11 1 2 3 9 9 9 9 9 9 19 9 
3 1 2 18 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 18 9 
6 1 2 3 20 19 9 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 18 21 16 
34 1 2 3 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 11 10 16 22 22 22 16 22 22 16 22 14 13 15 12 22 
3 1 2 18 
3 1 2 18 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
16 1 2 3 20 9 9 4 6 5 7 8 9 10 19 17 10 
19 1 2 3 20 4 5 6 7 8 9 10 11 10 16 13 14 12 15 16 
3 1 2 18 
20 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 11 10 18 21 16 
3 1 2 18 
22 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 11 10 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 19 17 
34 1 2 3 9 4 6 5 7 8 9 10 11 10 17 5 7 8 16 22 22 22 22 22 11 22 16 16 16 16 14 13 12 15 16 
14 1 2 3 4 5 6 7 8 9 10 10 10 19 17 
5 1 2 20 18 20 
4 1 2 18 20 
9 1 2 3 9 9 9 9 19 9 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
3 1 2 18 
32 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 16 16 16 16 16 16 18 21 16 
25 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 16 16 14 13 12 15 16 
19 1 2 3 20 9 9 9 4 5 6 7 8 9 10 11 10 21 18 16 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 20 9 19 9 
26 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 5 17 7 8 10 10 10 19 17 10 
3 1 2 18 
29 1 2 3 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 22 13 14 15 12 16 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 14 13 12 15 16 
21 1 2 3 20 9 9 4 5 6 7 8 9 11 10 16 16 14 12 15 13 16 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 13 14 12 15 16 
9 1 2 3 20 9 9 9 18 9 
15 1 2 3 20 4 6 5 7 8 9 10 10 10 19 17 
23 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
18 1 2 3 4 6 5 7 8 9 11 10 16 22 14 15 12 13 16 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 19 17 10 
21 1 2 20 3 20 9 4 6 5 7 8 9 10 10 10 11 10 16 18 21 22 
5 1 2 20 18 20 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
21 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 21 18 16 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 13 12 15 16 
3 1 2 18 
19 1 2 3 9 4 5 6 7 8 9 11 10 16 22 16 16 21 18 16 
27 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 16 16 16 16 16 16 13 14 12 15 16 
24 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 10 
18 1 2 3 9 4 9 5 6 7 8 9 11 10 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
6 1 2 3 9 19 9 
22 1 2 20 20 20 3 20 9 9 4 6 5 7 8 9 10 10 10 10 17 19 10 
27 1 2 3 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 14 15 13 12 16 
17 1 2 3 9 9 4 5 6 7 8 9 10 11 10 18 21 16 
6 1 2 3 9 18 9 
33 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 22 22 5 17 7 8 22 22 22 22 11 22 16 14 13 12 15 16 
3 1 2 18 
13 1 2 3 4 6 5 7 8 9 10 17 19 10 
56 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 10 10 10 10 10 10 10 10 10 10 10 10 
3 1 2 18 
18 1 2 3 20 4 6 5 7 8 9 5 17 7 8 10 17 19 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
23 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 17 19 
7 1 2 20 3 20 18 9 
15 1 2 3 9 4 5 6 7 8 9 11 10 16 19 17 
23 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
22 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 19 17 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
25 1 2 3 20 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 13 12 14 15 22 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
19 1 2 3 9 9 9 4 6 5 7 8 9 11 10 14 12 13 15 16 
31 1 2 20 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 16 16 16 13 14 12 15 16 
24 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 14 13 12 15 16 
24 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
18 1 2 3 20 4 6 5 7 8 9 10 11 10 14 12 13 15 16 
30 1 2 3 20 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 12 15 13 14 16 
14 1 2 3 20 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
5 1 2 3 18 9 
4 1 2 18 20 
3 1 2 18 
26 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 5 17 7 8 16 22 22 18 21 22 
31 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 22 16 16 22 22 14 13 12 15 16 
10 1 2 3 20 9 9 9 9 18 9 
5 1 2 3 19 9 
4 1 2 18 20 
26 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
17 1 2 3 9 4 5 6 7 8 9 11 10 13 15 14 12 16 
4 1 2 18 20 
5 1 2 3 18 9 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 10 10 21 18 10 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
24 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 14 15 13 12 16 
6 1 2 3 9 19 9 
10 1 2 3 9 9 9 9 9 9 19 
4 1 2 18 20 
15 1 2 3 9 4 5 6 7 8 9 10 10 19 17 10 
6 1 2 3 9 18 9 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 21 18 16 
25 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
14 1 2 3 4 6 5 7 8 9 10 10 10 17 19 
25 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 11 10 21 18 16 
25 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 15 14 12 13 16 
15 1 2 3 4 6 5 7 8 9 10 11 10 21 18 16 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 12 13 14 15 16 
3 1 2 18 
84 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 16 16 16 16 16 16 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 12 13 15 14 16 
4 1 2 18 20 
3 1 2 18 
9 1 2 3 9 9 9 9 19 9 
3 1 2 18 
15 1 2 3 9 4 6 5 7 8 9 11 10 21 18 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
19 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 
3 1 2 18 
9 1 2 3 9 9 9 9 18 9 
5 1 2 20 18 20 
21 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 18 21 16 
7 1 2 3 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
23 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 19 17 10 
3 1 2 18 
5 1 2 23 18 23 
44 1 2 3 9 9 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 14 13 12 15 16 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 9 9 4 6 5 7 8 9 11 10 16 22 22 18 21 22 
29 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 16 13 12 14 15 16 
27 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
26 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 14 12 13 15 16 
5 1 2 3 19 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 18 21 16 
3 1 2 18 
26 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 14 13 12 15 16 
4 1 2 18 20 
20 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 16 16 21 18 22 
14 1 2 3 4 5 6 7 8 9 10 10 10 17 19 
31 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 14 12 13 15 16 
27 1 2 3 9 4 5 6 7 8 9 11 10 17 5 7 8 16 22 22 22 11 22 14 12 13 15 16 
34 1 2 3 4 6 5 7 8 9 10 10 5 17 7 8 10 10 10 10 10 11 10 16 16 22 22 22 16 16 22 22 18 21 16 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
6 1 2 3 20 19 9 
3 1 2 18 
34 1 2 3 4 5 6 7 8 9 11 10 16 16 16 22 22 22 22 22 17 5 7 8 22 22 22 22 22 22 22 22 17 19 22 
12 1 2 3 4 6 5 7 8 9 19 17 10 
21 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 16 14 13 12 15 16 
5 1 2 3 18 9 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 14 13 15 12 16 
5 1 2 3 19 9 
15 1 2 3 9 4 5 6 7 8 9 10 10 10 17 19 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 11 10 16 21 18 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
46 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 11 10 5 17 7 8 16 22 22 22 22 11 22 13 14 15 12 16 
28 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 16 16 14 12 13 15 16 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 13 14 12 15 16 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
3 1 2 18 
19 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
25 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 5 17 7 8 10 11 10 21 18 16 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 11 10 18 21 16 
4 1 2 18 20 
15 1 2 3 9 9 4 6 5 7 8 9 10 21 18 10 
7 1 2 3 20 9 18 9 
18 1 2 3 20 4 6 5 7 8 9 10 11 10 13 14 15 12 16 
6 1 2 3 20 18 9 
3 1 2 18 
22 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 13 12 14 15 16 
3 1 2 18 
37 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 16 22 22 22 5 17 7 8 22 22 22 22 11 22 14 12 15 13 16 
21 1 2 3 4 6 5 7 8 9 11 10 16 16 22 22 22 14 12 13 15 16 
7 1 2 20 3 20 18 9 
4 1 2 18 20 
22 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 19 17 10 
26 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 22 22 14 12 13 15 16 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 11 10 16 16 19 17 16 
34 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 5 17 7 8 16 22 22 11 22 15 12 14 13 16 
51 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 19 17 10 
19 1 2 3 9 9 4 5 6 7 8 9 10 11 10 14 13 12 15 16 
3 1 2 18 
50 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 17 5 7 8 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 19 17 
17 1 2 3 9 4 6 5 7 8 9 10 11 10 16 18 21 16 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 14 12 13 15 16 
3 1 2 18 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 19 9 
4 1 2 18 20 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 13 12 15 16 
23 1 2 3 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 19 17 10 
16 1 2 3 4 5 6 7 8 9 11 10 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
31 1 2 3 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 17 5 7 8 10 10 11 10 14 13 12 15 16 
3 1 2 18 
47 1 2 3 20 9 9 4 9 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 11 10 16 17 5 7 8 16 13 14 12 15 22 
4 1 2 18 20 
8 1 2 3 20 9 9 19 9 
20 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
7 1 2 3 9 9 18 9 
3 1 2 18 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 11 10 16 16 22 22 22 13 15 12 14 16 
35 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 16 22 22 21 18 16 
26 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 16 16 14 13 15 12 16 
3 1 2 18 
5 1 2 20 18 20 
7 1 2 3 9 9 19 9 
7 1 2 3 4 9 19 9 
4 1 2 18 20 
3 1 2 18 
28 1 2 3 9 9 4 5 6 7 8 9 11 10 16 16 22 22 22 22 22 16 16 22 14 13 15 12 16 
10 1 2 3 20 9 9 9 9 18 9 
4 1 2 18 20 
20 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 13 14 12 15 16 
42 1 2 3 4 9 5 6 7 8 9 5 17 7 8 10 10 5 17 7 8 10 17 5 7 8 10 10 10 11 10 16 16 16 22 22 22 22 22 22 18 21 22 
39 1 2 3 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 16 16 22 22 22 22 16 16 13 14 15 12 16 
6 1 2 3 9 18 9 
17 1 2 20 20 3 20 4 6 5 7 8 9 10 10 17 19 10 
24 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 14 15 13 12 16 
3 1 2 18 
24 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
17 1 2 3 4 5 6 7 8 9 10 11 10 13 14 12 15 16 
5 1 2 3 18 9 
29 1 2 3 20 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
20 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 16 16 21 18 16 
6 1 2 3 4 19 9 
19 1 2 3 4 6 5 7 8 9 10 10 10 11 10 14 12 13 15 16 
27 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 14 12 15 13 22 
4 1 2 18 20 
4 1 2 18 20 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
26 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 17 5 7 8 16 14 15 13 12 22 
35 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 16 22 22 22 22 22 16 16 15 13 14 12 16 
66 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 9 18 9 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 12 13 15 14 16 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 10 10 11 10 21 18 16 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
22 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
14 1 2 3 9 9 4 5 6 7 8 9 17 19 10 
3 1 2 18 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 18 9 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
9 1 2 3 20 9 9 9 9 19 
22 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
18 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 19 17 10 
8 1 2 3 9 9 9 18 9 
3 1 2 18 
6 1 2 3 20 19 9 
3 1 2 18 
3 1 2 18 
28 1 2 3 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
4 1 2 18 20 
24 1 2 3 9 4 6 5 7 8 9 10 5 17 7 8 10 10 11 10 14 13 15 12 16 
18 1 2 3 9 4 5 6 7 8 9 11 10 16 14 13 15 12 16 
29 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 22 19 17 22 
36 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 17 5 7 8 10 10 11 10 16 22 22 22 22 16 16 14 13 12 15 16 
21 1 2 3 9 4 5 6 7 8 9 10 10 5 17 7 8 10 10 19 17 10 
3 1 2 18 
39 1 2 3 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
18 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
24 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 11 10 14 15 13 12 16 
5 1 2 3 19 9 
4 1 2 18 20 
3 1 2 18 
63 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 17 5 7 8 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 16 16 22 22 22 22 16 22 22 22 22 22 22 22 22 22 16 14 12 13 15 16 
17 1 2 3 9 9 4 6 5 7 8 9 10 11 10 18 21 16 
3 1 2 18 
22 1 2 3 9 9 4 5 6 7 8 9 11 10 16 22 22 22 14 13 15 12 16 
20 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 14 13 15 12 16 
4 1 2 18 20 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 9 19 
22 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 14 15 13 12 16 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 16 21 18 16 
42 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 17 5 7 8 10 10 10 11 10 16 22 22 22 16 22 22 22 22 22 22 22 14 13 15 12 16 
7 1 2 20 3 20 18 9 
5 1 2 20 18 20 
17 1 2 3 9 9 9 4 5 6 7 8 9 10 10 19 17 10 
9 1 2 20 20 20 20 20 18 20 
3 1 2 18 
57 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 14 13 15 12 16 
16 1 2 20 3 20 4 6 5 7 8 9 10 10 17 19 10 
3 1 2 18 
7 1 2 20 3 20 18 9 
4 1 2 18 20 
40 1 2 3 20 9 9 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
30 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 16 22 22 22 22 22 22 22 22 16 17 19 22 
25 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
21 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 10 17 19 10 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
33 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 14 12 13 15 16 
21 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 16 14 13 12 15 16 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
3 1 2 18 
59 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 17 5 7 8 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 13 14 12 15 16 
23 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 14 12 13 15 16 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
11 1 2 3 20 9 9 9 9 9 18 9 
22 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 12 14 13 15 16 
6 1 2 3 4 19 9 
32 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 22 22 16 17 5 7 8 16 14 12 13 15 22 
3 1 2 18 
21 1 2 3 20 9 9 4 5 6 7 8 9 10 10 11 10 13 14 15 12 16 
24 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 19 17 10 
20 1 2 3 9 9 9 4 9 6 5 7 8 9 11 10 13 12 14 15 16 
39 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
3 1 2 18 
19 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 
7 1 2 3 20 9 18 9 
28 1 2 3 20 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 21 18 16 
4 1 2 18 20 
6 1 2 3 20 18 9 
3 1 2 18 
18 1 2 3 9 9 4 5 6 7 8 9 11 10 14 15 13 12 16 
3 1 2 18 
24 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
10 1 2 3 9 9 9 9 9 9 19 
3 1 2 18 
14 1 2 3 9 9 4 5 6 7 8 9 19 17 10 
9 1 2 3 9 9 9 9 9 19 
11 1 2 23 23 20 23 20 20 20 18 20 
4 1 2 18 20 
16 1 2 3 4 6 5 7 8 9 10 10 11 10 18 21 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
13 1 2 3 9 4 5 6 7 8 9 17 19 10 
20 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 14 15 12 13 16 
3 1 2 18 
39 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 5 17 7 8 10 10 5 17 7 8 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
19 1 2 3 9 9 4 6 5 7 8 9 11 10 16 13 14 12 15 16 
3 1 2 18 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
22 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 11 10 14 13 12 15 16 
27 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
14 1 2 3 20 9 4 6 5 7 8 9 19 17 10 
12 1 2 3 4 5 6 7 8 9 19 17 10 
31 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
24 1 2 3 9 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 12 13 14 15 16 
43 1 2 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 17 5 7 8 16 15 13 14 12 22 
19 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
20 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 15 13 12 14 16 
22 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 21 18 16 
16 1 2 3 4 5 6 7 8 9 11 10 14 15 13 12 16 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
15 1 2 3 20 9 4 6 5 7 8 9 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
5 1 2 3 19 9 
23 1 2 3 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 21 18 16 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
23 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 16 16 12 13 14 15 16 
16 1 2 3 4 6 5 7 8 9 11 10 13 14 12 15 16 
5 1 2 20 18 20 
6 1 2 20 20 18 20 
24 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 16 22 13 14 15 12 16 
6 1 2 23 23 18 23 
3 1 2 18 
6 1 2 20 20 18 20 
3 1 2 18 
3 1 2 18 
26 1 2 20 20 20 20 20 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 10 17 19 10 
18 1 2 20 20 3 20 4 6 5 7 8 9 10 10 10 21 18 10 
4 1 2 18 20 
3 1 2 18 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
7 1 2 20 3 20 18 9 
24 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 14 15 13 12 16 
53 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 16 14 12 13 15 16 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 17 19 22 
27 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 10 11 10 13 15 12 14 16 
5 1 2 20 18 20 
5 1 2 20 18 20 
24 1 2 3 20 4 9 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 10 19 17 
3 1 2 18 
22 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 18 21 16 
5 1 2 20 18 20 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
5 1 2 3 19 9 
19 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 19 17 
25 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
20 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
19 1 2 3 9 9 4 6 5 7 8 9 10 11 10 12 14 15 13 16 
19 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
5 1 2 20 18 20 
3 1 2 18 
31 1 2 3 4 9 5 6 7 8 9 10 5 17 7 8 10 11 10 16 16 16 5 17 7 8 16 13 14 12 15 22 
25 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 11 10 13 14 15 12 16 
7 1 2 3 20 9 18 9 
34 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 16 16 16 17 5 7 8 16 14 15 13 12 22 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 12 13 15 16 
4 1 2 18 20 
27 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
9 1 2 3 9 9 9 9 19 9 
15 1 2 3 4 5 6 7 8 9 10 10 10 19 17 10 
7 1 2 3 9 9 19 9 
32 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 22 17 5 7 8 16 13 14 12 15 22 
3 1 2 18 
4 1 2 18 20 
38 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 17 19 
28 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 19 17 
21 1 2 3 4 9 5 6 7 8 9 10 10 10 10 11 10 14 13 15 12 16 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 17 19 10 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 19 17 10 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 11 10 14 12 13 15 16 
21 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 14 13 15 12 22 
3 1 2 18 
15 1 2 3 9 4 5 6 7 8 9 10 10 19 17 10 
24 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 21 18 16 
5 1 2 20 18 20 
4 1 2 18 20 
10 1 2 3 9 9 9 9 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 9 9 19 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
69 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 12 15 13 14 16 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
36 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 21 18 16 
3 1 2 18 
6 1 2 3 9 18 9 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 21 18 10 
4 1 2 18 20 
13 1 2 3 20 4 5 6 7 8 9 19 17 10 
22 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 19 17 10 
5 1 2 20 18 20 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
16 1 2 3 20 4 5 6 7 8 9 10 10 10 17 19 10 
22 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 11 10 16 16 21 18 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
22 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 19 17 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
7 1 2 3 20 9 18 9 
6 1 2 3 20 19 9 
31 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 11 10 21 18 16 
16 1 2 3 4 5 6 7 8 9 11 10 14 12 13 15 16 
3 1 2 18 
29 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 16 16 16 14 15 13 12 16 
28 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 16 22 22 22 12 13 15 14 16 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
6 1 2 20 20 18 20 
4 1 2 18 20 
5 1 2 20 18 20 
3 1 2 18 
5 1 2 3 19 9 
19 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 18 21 16 
26 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 22 22 22 22 22 22 22 17 19 22 
18 1 2 3 9 9 4 5 6 7 8 9 11 10 13 14 15 12 16 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 19 9 
4 1 2 18 20 
16 1 2 3 20 9 4 5 6 7 8 9 10 10 17 19 10 
35 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 17 5 7 8 10 10 11 10 16 22 22 22 22 16 14 13 15 12 16 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 10 17 19 
22 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 18 21 16 
24 1 2 20 3 20 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 18 21 22 
25 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 19 17 10 
3 1 2 18 
33 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 11 10 16 16 16 22 22 22 22 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
23 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 16 16 16 16 18 21 22 
4 1 2 18 20 
85 1 2 3 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 16 16 16 16 16 16 16 16 16 16 16 16 16 16 16 16 16 16 16 16 16 16 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 16 22 22 22 22 22 22 22 22 19 17 22 
3 1 2 18 
33 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 18 9 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 13 15 12 14 16 
3 1 2 18 
26 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 16 14 12 13 15 16 
15 1 2 3 4 6 5 7 8 9 10 10 10 19 17 10 
19 1 2 3 4 6 5 7 8 9 10 11 10 16 16 12 14 13 15 16 
28 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 15 13 12 14 16 
37 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 17 5 7 8 10 10 17 5 7 8 10 10 10 11 10 16 18 21 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
14 1 2 20 3 20 9 9 9 9 9 9 9 18 9 
24 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 16 22 19 17 22 
19 1 2 3 20 4 6 5 7 8 9 10 11 10 16 14 13 15 12 16 
29 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 14 15 13 12 16 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 14 15 13 12 16 
4 1 2 18 20 
32 1 2 3 9 9 4 6 5 7 8 9 10 10 10 17 5 7 8 10 10 10 10 11 10 16 22 22 16 22 19 17 22 
22 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 16 22 22 21 18 22 
26 1 2 3 9 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 17 19 10 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 19 17 10 
22 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 11 10 13 14 12 15 16 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 21 18 16 
27 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
19 1 2 3 9 4 6 5 7 8 9 10 10 11 10 13 15 14 12 16 
20 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 17 19 10 
25 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 16 16 16 16 14 15 12 13 16 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
18 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
29 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 13 12 14 15 16 
6 1 2 3 20 19 9 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 18 21 16 
24 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 14 12 15 13 16 
3 1 2 18 
8 1 2 20 20 3 20 18 9 
20 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 13 14 12 15 16 
17 1 2 3 4 5 6 7 8 9 10 11 10 12 13 15 14 16 
5 1 2 3 19 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
19 1 2 3 20 4 6 5 7 8 9 10 11 10 16 14 13 15 12 16 
3 1 2 18 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 9 9 19 9 
26 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 5 17 7 8 10 11 10 18 21 16 
3 1 2 18 
29 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 11 10 18 21 16 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
73 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
21 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 12 13 15 14 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
11 1 2 20 3 20 9 9 9 9 18 9 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 10 10 11 10 12 15 14 13 16 
6 1 2 3 9 19 9 
16 1 2 3 4 5 6 7 8 9 11 10 14 15 13 12 16 
6 1 2 3 20 19 9 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
13 1 2 3 4 6 5 7 8 9 10 17 19 10 
27 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 16 14 12 13 15 16 
7 1 2 3 9 9 18 9 
6 1 2 3 20 18 9 
4 1 2 18 20 
70 1 2 3 20 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 16 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 22 11 22 16 22 22 22 22 22 22 22 22 16 13 14 15 12 16 
20 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 19 17 
4 1 2 18 20 
4 1 2 18 20 
25 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 16 22 22 22 22 13 14 15 12 16 
20 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 14 13 12 15 16 
59 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 5 17 7 8 10 10 10 11 10 17 5 7 8 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 13 14 15 12 16 
3 1 2 18 
62 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 5 17 7 8 10 17 5 7 8 10 10 10 11 10 16 22 5 17 7 8 22 22 5 17 7 8 22 22 5 17 7 8 22 22 22 22 22 22 22 11 22 13 14 15 12 16 
4 1 2 18 20 
4 1 2 18 20 
20 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 14 12 13 15 16 
13 1 2 3 9 4 6 5 7 8 9 17 19 10 
46 1 2 3 20 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 16 16 16 22 22 22 22 16 22 22 22 22 22 22 22 22 22 14 13 12 15 16 
7 1 2 20 20 20 18 20 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 17 19 10 
8 1 2 20 3 20 9 18 9 
19 1 2 3 20 4 6 5 7 8 9 10 10 10 10 11 10 21 18 16 
6 1 2 3 20 18 9 
30 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 16 16 16 15 12 14 13 16 
25 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
31 1 2 3 4 9 6 5 7 8 9 5 17 7 8 10 10 5 17 7 8 10 10 11 10 16 22 16 16 18 21 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
23 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 15 14 13 12 16 
31 1 2 3 9 4 6 5 7 8 9 10 11 10 16 5 17 7 8 16 22 22 22 22 22 11 22 14 12 13 15 16 
5 1 2 3 19 9 
30 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
8 1 2 3 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
24 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 13 14 15 12 16 
7 1 2 3 9 9 18 9 
10 1 2 3 9 9 9 9 9 19 9 
29 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
27 1 2 3 9 4 5 6 7 8 9 11 10 16 16 16 22 22 16 22 22 22 22 13 12 14 15 16 
4 1 2 18 20 
17 1 2 3 4 5 6 7 8 9 10 11 10 16 16 18 21 16 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
39 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 22 16 22 22 22 22 16 22 22 15 12 14 13 16 
28 1 2 3 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 16 14 13 12 15 16 
3 1 2 18 
24 1 2 3 20 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 19 17 10 
36 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 11 10 16 16 16 14 13 15 12 16 
8 1 2 3 20 9 9 18 9 
5 1 2 20 18 20 
6 1 2 3 9 19 9 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 20 9 18 9 
21 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 14 12 13 15 16 
6 1 2 3 20 18 9 
3 1 2 18 
6 1 2 20 20 18 20 
19 1 2 20 3 20 9 9 9 9 4 6 5 7 8 9 10 19 17 10 
3 1 2 18 
6 1 2 3 20 18 9 
29 1 2 3 4 5 6 7 8 9 17 5 7 8 10 11 10 16 22 22 16 16 22 22 22 13 12 15 14 16 
14 1 2 3 4 5 6 7 8 9 10 10 17 19 10 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 19 9 
7 1 2 3 20 9 19 9 
3 1 2 18 
7 1 2 3 9 9 19 9 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 14 12 13 15 16 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 18 21 16 
16 1 2 20 3 20 9 4 5 6 7 8 9 10 19 17 10 
4 1 2 18 20 
6 1 2 3 9 18 9 
12 1 2 3 4 6 5 7 8 9 17 19 10 
33 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 16 22 22 22 16 16 16 16 16 22 22 22 16 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
26 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 14 15 13 12 16 
17 1 2 3 4 5 6 7 8 9 10 11 10 15 13 12 14 16 
16 1 2 3 4 5 6 7 8 9 11 10 14 13 12 15 16 
5 1 2 20 18 20 
3 1 2 18 
12 1 2 3 20 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 19 9 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
6 1 2 20 20 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 11 10 14 15 13 12 16 
6 1 2 3 20 18 9 
22 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 18 21 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 20 18 20 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 20 4 5 6 7 8 9 11 10 16 14 12 15 13 16 
3 1 2 18 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 10 11 10 16 14 13 12 15 16 
11 1 2 3 20 9 9 9 9 9 18 9 
3 1 2 18 
19 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 16 18 21 16 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 3 18 9 
3 1 2 18 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 18 21 16 
3 1 2 18 
38 1 2 3 9 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
42 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 16 22 22 16 16 22 22 22 22 22 22 22 22 16 16 16 16 14 15 13 12 16 
10 1 2 3 9 9 9 9 9 18 9 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
6 1 2 3 9 19 9 
4 1 2 18 20 
7 1 2 23 23 23 18 23 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 9 18 9 
20 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 13 14 12 15 16 
10 1 2 3 9 9 9 9 9 18 9 
38 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 17 5 7 8 10 10 10 10 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 11 10 16 22 22 14 12 15 13 16 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
40 1 2 3 20 4 6 5 7 8 9 10 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 17 5 7 8 22 22 22 11 22 13 14 12 15 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
27 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 14 13 12 15 16 
7 1 2 3 9 9 18 9 
3 1 2 18 
9 1 2 20 20 20 20 20 18 20 
4 1 2 18 20 
24 1 2 20 20 20 20 20 20 20 3 20 4 5 6 7 8 9 11 10 13 14 15 12 16 
5 1 2 20 18 20 
5 1 2 20 18 20 
5 1 2 20 18 20 
13 1 2 3 20 4 5 6 7 8 9 17 19 10 
4 1 2 18 20 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
6 1 2 3 20 19 9 
6 1 2 20 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
20 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 17 19 10 
4 1 2 18 20 
18 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
26 1 2 20 20 20 20 20 3 20 4 6 5 7 8 9 10 10 10 10 11 10 12 13 15 14 16 
6 1 2 20 23 18 23 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
34 1 2 3 20 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 11 10 16 22 22 22 16 22 22 22 15 12 13 14 16 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
30 1 2 20 3 20 9 9 4 6 5 7 8 9 5 17 7 8 10 11 10 17 5 7 8 16 14 12 15 13 22 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
26 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 16 18 21 22 
17 1 2 3 9 9 4 6 5 7 8 9 10 10 10 19 17 10 
6 1 2 3 9 18 9 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 18 9 
11 1 2 3 20 9 9 9 9 9 18 9 
9 1 2 3 9 9 9 9 18 9 
6 1 2 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 17 19 10 
7 1 2 3 20 9 18 9 
33 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
32 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 17 5 7 8 10 10 10 11 10 16 14 15 12 13 16 
19 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
28 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 16 16 22 22 14 12 15 13 16 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
11 1 2 3 9 9 9 9 9 9 19 9 
3 1 2 18 
26 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
28 1 2 3 20 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 21 18 16 
35 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 19 9 
23 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 16 15 13 14 12 16 
25 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 14 12 15 13 16 
3 1 2 18 
3 1 2 18 
5 1 2 3 18 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
14 1 2 3 9 4 5 6 7 8 9 10 18 21 10 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
6 1 2 20 20 18 20 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 20 18 20 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
6 1 2 3 20 18 9 
5 1 2 20 18 20 
22 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
16 1 2 3 4 5 6 7 8 9 10 10 11 10 21 18 16 
3 1 2 18 
26 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 11 10 13 14 15 12 16 
5 1 2 3 19 9 
35 1 2 3 4 6 5 7 8 9 17 5 7 8 10 5 17 7 8 10 10 5 17 7 8 10 10 10 10 11 10 14 13 15 12 16 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 9 19 9 
19 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 17 19 10 
26 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 16 16 16 14 13 12 15 16 
26 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 16 13 14 12 15 16 
3 1 2 18 
30 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 20 9 18 9 
5 1 2 3 19 9 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
4 1 2 18 20 
5 1 2 20 18 20 
23 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 11 10 14 13 12 15 16 
34 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 17 5 7 8 10 10 11 10 16 22 22 22 22 22 22 21 18 16 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
23 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 16 22 22 12 15 13 14 16 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
10 1 2 3 20 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 12 13 15 14 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
17 1 2 3 9 9 4 5 6 7 8 9 11 10 16 18 21 16 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
25 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 12 14 13 15 16 
3 1 2 18 
3 1 2 18 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
10 1 2 3 20 9 9 9 9 19 9 
17 1 2 3 20 9 4 6 5 7 8 9 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
5 1 2 23 18 23 
15 1 2 3 9 9 9 4 6 5 7 8 9 19 17 10 
24 1 2 3 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 14 12 13 15 16 
38 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 11 10 16 22 22 22 16 22 22 22 22 14 13 12 15 16 
30 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 17 5 7 8 16 12 14 15 13 22 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
18 1 2 3 20 9 4 6 5 7 8 9 11 10 14 12 13 15 16 
11 1 2 20 20 20 20 20 20 20 18 20 
16 1 2 3 9 4 6 5 7 8 9 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
13 1 2 3 4 6 5 7 8 9 10 17 19 10 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 9 9 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
21 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
58 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 16 
24 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 16 22 22 13 14 12 15 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
23 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 14 13 15 12 16 
3 1 2 18 
22 1 2 20 3 20 4 5 6 7 8 9 10 11 10 16 16 22 13 15 12 14 16 
15 1 2 3 9 4 6 5 7 8 9 11 10 18 21 16 
10 1 2 3 9 9 9 9 9 19 9 
3 1 2 18 
6 1 2 3 20 18 9 
5 1 2 3 19 9 
41 1 2 3 9 9 9 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 14 13 12 15 16 
7 1 2 3 20 9 18 9 
12 1 2 3 9 9 9 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
31 1 2 3 20 9 9 4 6 5 7 8 9 5 17 7 8 10 17 5 7 8 10 10 10 11 10 13 14 15 12 16 
5 1 2 20 18 20 
22 1 2 3 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 19 17 10 
4 1 2 18 20 
5 1 2 23 18 23 
3 1 2 18 
20 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 10 17 19 10 
4 1 2 18 20 
5 1 2 3 18 9 
11 1 2 3 9 9 9 9 9 9 19 9 
38 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 16 16 17 5 7 8 16 22 22 22 22 11 22 14 12 13 15 16 
20 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 14 12 13 15 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
25 1 2 3 9 4 6 5 7 8 9 10 5 17 7 8 10 10 11 10 16 14 13 15 12 16 
8 1 2 3 20 9 9 18 9 
21 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
16 1 2 3 4 6 5 7 8 9 11 10 13 14 12 15 16 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
20 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 11 10 21 18 16 
24 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 14 15 12 13 16 
40 1 2 3 20 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 10 10 5 17 7 8 10 10 10 10 11 10 16 16 22 22 14 13 12 15 22 
48 1 2 3 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 11 10 10 10 10 10 14 12 13 15 16 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
21 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 18 21 16 
9 1 2 3 20 9 9 9 18 9 
21 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 16 14 12 13 15 16 
6 1 2 3 20 18 9 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 18 21 16 
4 1 2 18 20 
37 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 11 10 14 12 13 15 16 
4 1 2 18 20 
21 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 14 13 12 15 16 
10 1 2 20 3 20 9 9 9 18 9 
33 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
24 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
29 1 2 3 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 11 10 14 12 13 15 16 
3 1 2 18 
25 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
7 1 2 3 20 9 18 9 
3 1 2 18 
20 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 19 17 
24 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 16 14 15 13 12 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
22 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 11 10 13 14 15 12 16 
6 1 2 3 9 19 9 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
14 1 2 3 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
14 1 2 3 9 9 4 6 5 7 8 9 17 19 10 
9 1 2 3 20 9 9 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
11 1 2 3 20 9 9 9 9 9 18 9 
3 1 2 18 
16 1 2 3 9 9 9 4 5 6 7 8 9 10 10 19 17 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
15 1 2 3 20 9 9 9 9 9 9 9 4 9 19 9 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 4 5 6 7 8 9 11 10 16 22 22 14 13 12 15 16 
33 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 16 16 22 22 16 16 16 14 13 15 12 16 
43 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 17 5 7 8 10 17 5 7 8 10 10 10 11 10 16 22 22 22 18 21 22 
4 1 2 18 20 
26 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 11 10 14 13 12 15 16 
3 1 2 18 
7 1 2 3 9 9 19 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
17 1 2 3 9 9 9 9 4 6 5 7 8 9 10 19 17 10 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
31 1 2 20 3 20 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 18 21 16 
4 1 2 18 20 
42 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 16 16 16 22 22 22 22 16 16 22 22 22 22 17 19 22 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
28 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
14 1 2 3 4 5 6 7 8 9 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 19 9 
6 1 2 3 20 18 9 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 14 15 12 13 16 
28 1 2 3 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
9 1 2 3 9 9 9 9 19 9 
3 1 2 18 
23 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 12 13 14 15 16 
3 1 2 18 
38 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 16 22 14 12 13 15 22 
15 1 2 3 9 4 5 6 7 8 9 10 10 19 17 10 
37 1 2 20 20 20 20 20 20 3 20 9 9 9 9 4 9 6 5 7 8 9 10 11 10 16 22 22 22 16 22 22 16 14 12 13 15 16 
3 1 2 18 
9 1 2 3 9 9 9 4 19 9 
17 1 2 3 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
36 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 16 16 16 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
17 1 2 3 9 4 5 6 7 8 9 10 10 11 10 18 21 16 
5 1 2 23 18 23 
8 1 2 3 9 9 9 18 9 
15 1 2 3 9 4 5 6 7 8 9 11 10 21 18 16 
3 1 2 18 
29 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 10 10 10 10 10 17 19 10 
22 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 11 10 14 13 12 15 16 
14 1 2 3 20 4 5 6 7 8 9 10 17 19 10 
3 1 2 18 
21 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
29 1 2 3 9 9 9 4 9 6 5 7 8 9 10 10 17 5 7 8 10 10 10 11 10 14 12 15 13 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 21 18 16 
5 1 2 3 18 9 
30 1 2 20 20 3 20 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 16 21 18 16 
4 1 2 18 20 
6 1 2 3 9 18 9 
4 1 2 18 20 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 14 12 15 13 16 
28 1 2 3 4 6 5 7 8 9 10 11 10 16 5 17 7 8 16 22 22 22 11 22 14 12 13 15 16 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
4 1 2 18 20 
16 1 2 3 20 9 4 6 5 7 8 9 10 10 19 17 10 
23 1 2 3 20 4 5 6 7 8 9 10 5 17 7 8 10 11 10 14 15 13 12 16 
4 1 2 18 20 
6 1 2 20 20 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 11 10 16 16 18 21 16 
12 1 2 3 20 9 9 9 9 9 9 18 9 
6 1 2 3 20 18 9 
7 1 2 3 20 9 19 9 
28 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 11 10 18 21 16 
30 1 2 3 9 9 4 6 5 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 10 10 11 10 18 21 16 
20 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 14 12 15 13 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 10 11 10 16 12 13 14 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 13 15 12 16 
5 1 2 23 18 23 
47 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 5 17 7 8 10 10 17 5 7 8 10 5 17 7 8 10 10 10 10 10 10 11 10 14 12 13 15 16 
4 1 2 18 20 
47 1 2 3 4 5 6 7 8 9 10 10 11 10 16 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 14 12 15 13 16 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 15 13 12 16 
42 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
4 1 2 18 20 
34 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 22 22 14 13 12 15 16 
5 1 2 3 18 9 
7 1 2 3 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
15 1 2 3 9 9 4 5 6 7 8 9 10 19 17 10 
20 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 12 15 13 14 16 
18 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 17 19 10 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 17 19 10 
17 1 2 3 9 4 6 5 7 8 9 10 10 10 10 19 17 10 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
24 1 2 3 20 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 10 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 9 19 9 
3 1 2 18 
4 1 2 18 20 
42 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 16 18 21 16 
26 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 16 16 18 21 16 
9 1 2 3 9 9 9 9 19 9 
4 1 2 18 20 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
12 1 2 3 9 9 9 9 9 9 9 19 9 
20 1 2 3 20 4 5 6 7 8 9 10 11 10 16 16 15 13 12 14 16 
15 1 2 3 9 4 6 5 7 8 9 11 10 18 21 16 
20 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 14 13 15 12 16 
5 1 2 20 18 20 
37 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 11 10 16 16 22 22 22 22 16 16 22 22 12 14 13 15 16 
4 1 2 18 20 
3 1 2 18 
29 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 16 15 12 13 14 16 
4 1 2 18 20 
37 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
11 1 2 3 20 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
22 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 22 22 14 12 13 15 16 
19 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 19 17 10 
22 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 22 22 14 13 12 15 16 
10 1 2 3 9 9 9 9 9 19 9 
16 1 2 3 4 6 5 7 8 9 11 10 12 13 15 14 16 
56 1 2 3 20 9 4 5 6 7 8 9 10 5 17 7 8 10 10 11 10 16 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 22 11 22 16 13 12 14 15 16 
26 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 19 17 10 
23 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 21 18 22 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 14 15 13 12 16 
4 1 2 18 20 
6 1 2 3 9 19 9 
23 1 2 3 20 4 5 6 7 8 9 10 11 10 16 16 22 22 22 12 14 13 15 16 
4 1 2 18 20 
9 1 2 3 9 9 9 9 19 9 
4 1 2 18 20 
5 1 2 3 19 9 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 9 18 9 
19 1 2 3 9 9 4 6 5 7 8 9 10 11 10 12 14 13 15 16 
7 1 2 3 20 9 18 9 
3 1 2 18 
23 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 22 16 12 14 13 15 16 
14 1 2 3 20 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
27 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 16 13 14 15 12 16 
5 1 2 20 18 20 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 18 9 
31 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
96 1 2 3 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 17 5 7 8 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 19 17 22 
3 1 2 18 
23 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 17 19 10 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 14 12 13 15 16 
14 1 2 3 4 5 6 7 8 9 11 10 18 21 16 
17 1 2 3 20 4 5 6 7 8 9 10 10 10 10 17 19 10 
4 1 2 18 20 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
17 1 2 3 20 9 4 6 5 7 8 9 10 10 10 17 19 10 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
8 1 2 3 9 9 9 18 9 
4 1 2 18 20 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
16 1 2 3 9 9 9 4 6 5 7 8 9 10 19 17 10 
29 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 16 22 22 16 14 15 13 12 16 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 17 19 16 
4 1 2 18 20 
10 1 2 3 9 9 9 9 9 18 9 
15 1 2 3 9 4 6 5 7 8 9 11 10 18 21 16 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
21 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
9 1 2 3 20 9 9 9 18 9 
24 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
28 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 19 17 10 
16 1 2 3 4 6 5 7 8 9 10 11 10 16 18 21 16 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 13 14 12 15 16 
18 1 2 3 20 4 5 6 7 8 9 10 11 10 12 14 13 15 16 
3 1 2 18 
25 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 16 14 13 12 15 16 
5 1 2 20 18 20 
3 1 2 18 
36 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 16 16 16 16 22 22 22 16 22 22 22 22 22 22 22 22 22 22 19 17 22 
4 1 2 18 20 
13 1 2 3 4 6 5 7 8 9 10 17 19 10 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 11 10 14 12 13 15 16 
4 1 2 18 20 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
31 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 14 12 15 13 16 
3 1 2 18 
25 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 13 14 15 12 16 
10 1 2 3 9 9 9 9 9 18 9 
18 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 17 19 10 
9 1 2 3 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 4 6 5 7 8 9 11 10 14 13 15 12 16 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 19 9 
12 1 2 3 9 9 9 9 9 9 9 19 9 
3 1 2 18 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
38 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 16 16 22 22 22 22 16 16 16 22 22 22 22 12 15 13 14 16 
33 1 2 3 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 11 10 16 16 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 16 16 21 18 16 
3 1 2 18 
36 1 2 3 4 6 5 7 8 9 10 11 10 16 23 16 16 22 22 22 22 22 22 22 22 22 22 22 22 16 16 22 13 14 15 12 16 
44 1 2 20 3 20 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 5 17 7 8 10 10 10 11 10 16 22 22 22 16 16 16 16 14 13 15 12 16 
4 1 2 18 20 
28 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
17 1 2 3 9 4 5 6 7 8 9 11 10 13 12 14 15 16 
5 1 2 3 19 9 
25 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 16 13 14 12 15 16 
21 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 17 19 22 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
38 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 5 17 7 8 16 22 22 22 22 22 22 22 22 22 22 22 11 22 14 12 13 15 16 
15 1 2 3 4 6 5 7 8 9 10 10 10 10 17 19 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
28 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 17 5 7 8 16 15 13 12 14 22 
4 1 2 18 20 
5 1 2 23 18 23 
4 1 2 18 20 
24 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 14 13 12 15 16 
6 1 2 3 9 18 9 
12 1 2 3 9 9 9 9 9 9 9 9 19 
5 1 2 20 18 20 
28 1 2 3 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 17 19 
9 1 2 3 20 9 9 9 19 9 
4 1 2 18 20 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
21 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 21 18 16 
6 1 2 3 20 18 9 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 12 14 13 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
18 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 3 18 9 
5 1 2 20 18 20 
4 1 2 18 20 
27 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 13 14 15 12 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
48 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 16 16 22 22 22 22 16 16 16 16 16 16 16 22 22 22 22 22 5 17 7 8 22 22 22 11 22 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 19 9 
3 1 2 18 
22 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 14 12 15 13 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 18 21 16 
3 1 2 18 
26 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 16 22 22 22 22 22 22 19 17 22 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 23 18 23 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 21 18 22 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
17 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 19 9 
34 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 22 16 14 15 13 12 16 
3 1 2 18 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
16 1 2 3 20 9 4 5 6 7 8 9 11 10 18 21 16 
5 1 2 20 18 20 
30 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 16 21 18 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 18 9 
6 1 2 3 9 18 9 
22 1 2 3 4 6 5 7 8 9 11 10 16 22 22 16 22 22 13 14 15 12 16 
24 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 16 16 22 22 14 13 12 15 16 
9 1 2 3 9 9 9 9 18 9 
3 1 2 18 
27 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 16 15 12 14 13 16 
26 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
5 1 2 20 18 20 
6 1 2 3 9 19 9 
41 1 2 3 9 4 6 5 7 8 9 10 5 17 7 8 10 10 17 5 7 8 10 5 17 7 8 10 10 11 10 16 16 16 16 22 22 22 22 19 17 22 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
20 1 2 20 3 20 9 4 5 6 7 8 9 11 10 16 14 13 12 15 16 
28 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 5 17 7 8 10 10 11 10 16 16 18 21 16 
3 1 2 18 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 12 15 13 16 
4 1 2 18 20 
5 1 2 3 19 9 
5 1 2 20 18 20 
24 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
23 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 3 19 9 
27 1 2 3 20 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 16 16 22 14 12 13 15 16 
35 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 16 16 16 16 22 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 13 12 14 15 16 
4 1 2 18 20 
15 1 2 3 9 9 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
11 1 2 20 3 20 9 9 9 9 19 9 
27 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 16 12 15 14 13 16 
5 1 2 20 18 20 
4 1 2 18 20 
36 1 2 3 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 16 5 17 7 8 22 22 22 11 22 14 15 12 13 16 
6 1 2 3 20 18 9 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
14 1 2 3 20 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
3 1 2 18 
25 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
7 1 2 20 20 20 18 20 
4 1 2 18 20 
27 1 2 20 20 20 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 14 12 13 15 16 
5 1 2 3 19 9 
22 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 13 14 12 15 16 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
42 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 15 12 14 13 16 
18 1 2 3 9 4 6 5 7 8 9 11 10 16 14 15 12 13 16 
3 1 2 18 
3 1 2 18 
28 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 5 17 7 8 10 10 11 10 18 21 16 
3 1 2 18 
34 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
32 1 2 3 4 6 5 7 8 9 10 10 10 10 10 11 10 16 16 16 16 16 22 22 22 22 22 22 13 14 12 15 16 
5 1 2 3 19 9 
7 1 2 3 9 9 19 9 
7 1 2 3 9 9 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
34 1 2 3 20 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 10 11 10 16 16 16 16 16 16 14 13 12 15 16 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
5 1 2 3 18 9 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 3 19 9 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
4 1 2 18 20 
7 1 2 20 3 20 18 9 
4 1 2 18 20 
27 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 20 18 9 
16 1 2 3 9 4 6 5 7 8 9 11 10 16 18 21 16 
13 1 2 3 20 9 9 9 9 9 9 9 9 19 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
30 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 22 21 18 16 
10 1 2 20 3 20 9 9 9 9 19 
26 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 16 16 14 12 15 13 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 17 19 10 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
9 1 2 3 20 9 9 9 19 9 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
18 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
16 1 2 3 20 4 5 6 7 8 9 10 10 10 19 17 10 
28 1 2 3 9 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 17 19 22 
19 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 19 17 10 
3 1 2 18 
24 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 17 19 22 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
23 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 9 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 18 21 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
39 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
25 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
5 1 2 23 18 23 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
6 1 2 3 9 18 9 
22 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 22 12 14 13 15 16 
27 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 20 18 20 
5 1 2 20 18 20 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 17 19 
5 1 2 20 18 20 
11 1 2 3 9 9 9 9 9 9 19 9 
7 1 2 3 9 9 18 9 
7 1 2 3 9 9 19 9 
7 1 2 20 3 20 18 9 
9 1 2 20 20 20 20 20 18 20 
7 1 2 3 9 9 18 9 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
30 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 16 16 22 22 22 22 22 22 22 12 14 13 15 16 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
13 1 2 3 9 4 6 5 7 8 9 17 19 10 
3 1 2 18 
48 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 5 17 7 8 10 10 10 11 10 16 16 23 16 16 22 22 22 22 22 22 22 22 16 16 14 13 15 12 16 
3 1 2 18 
21 1 2 3 9 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 19 17 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
20 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 13 12 14 15 16 
5 1 2 20 18 20 
9 1 2 3 20 9 9 9 18 9 
6 1 2 3 20 18 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
26 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
15 1 2 3 20 4 6 5 7 8 9 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 20 18 9 
26 1 2 3 9 9 4 6 5 7 8 9 10 10 17 5 7 8 10 10 11 10 14 15 13 12 16 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 20 4 6 5 7 8 9 11 10 14 12 13 15 16 
3 1 2 18 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
6 1 2 3 9 19 9 
6 1 2 3 20 18 9 
3 1 2 18 
4 1 2 18 20 
33 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
9 1 2 3 20 9 9 9 19 9 
3 1 2 18 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
6 1 2 3 4 19 9 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 11 10 16 14 12 13 15 16 
5 1 2 3 18 9 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
25 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 14 13 12 15 16 
5 1 2 3 19 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 20 18 20 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
5 1 2 23 18 23 
46 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 16 22 22 22 22 22 22 14 12 13 15 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 19 17 10 
4 1 2 18 20 
5 1 2 20 18 20 
20 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 13 14 12 15 16 
5 1 2 20 18 20 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 21 18 16 
4 1 2 18 20 
3 1 2 18 
26 1 2 3 20 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
19 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
3 1 2 18 
22 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 21 18 16 
16 1 2 3 20 4 5 6 7 8 9 10 10 10 19 17 10 
22 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 13 14 12 15 16 
21 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 18 21 22 
24 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
34 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
24 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
14 1 2 20 3 20 4 6 5 7 8 9 19 17 10 
4 1 2 18 20 
6 1 2 3 20 18 9 
9 1 2 3 20 9 9 9 18 9 
61 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 5 17 7 8 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 16 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 19 17 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
23 1 2 3 9 9 4 6 5 7 8 9 11 10 16 22 22 16 16 14 13 12 15 16 
9 1 2 3 9 9 9 9 19 9 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 16 21 18 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
28 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 15 13 12 14 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
9 1 2 20 20 3 20 9 18 9 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 19 9 
29 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 16 16 22 22 22 12 13 15 14 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
23 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
7 1 2 3 20 9 9 19 
20 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 17 19 10 
65 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 10 17 5 7 8 10 5 17 7 8 10 5 17 7 8 10 5 17 7 8 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 5 17 7 8 16 14 12 13 15 22 
3 1 2 18 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
24 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 18 21 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
15 1 2 3 4 5 6 7 8 9 10 11 10 18 21 16 
71 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 22 22 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
4 1 2 18 20 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
26 1 2 20 20 20 20 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 18 21 16 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
6 1 2 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
29 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 14 13 15 12 16 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 18 9 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 11 10 16 16 12 14 15 13 16 
33 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 16 22 22 22 22 22 22 14 13 12 15 16 
4 1 2 18 20 
33 1 2 20 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 22 17 5 7 8 22 22 22 11 22 14 12 15 13 16 
4 1 2 18 20 
34 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 5 17 7 8 10 10 10 10 10 10 10 11 10 16 14 13 12 15 16 
3 1 2 18 
35 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 11 10 16 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 10 10 10 10 11 10 16 14 13 12 15 16 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 20 18 9 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 14 15 12 13 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
6 1 2 3 20 18 9 
6 1 2 3 20 18 9 
6 1 2 3 9 18 9 
17 1 2 3 9 4 6 5 7 8 9 11 10 12 14 15 13 16 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 14 13 12 15 16 
3 1 2 18 
39 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 11 10 17 5 7 8 16 22 22 22 22 22 22 22 22 22 22 11 22 14 13 15 12 16 
18 1 2 3 4 5 6 7 8 9 11 10 16 16 15 12 14 13 16 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 13 15 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
26 1 2 3 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 11 10 16 21 18 16 
7 1 2 3 9 9 19 9 
3 1 2 18 
35 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 5 17 7 8 10 10 19 17 10 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
3 1 2 18 
28 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
42 1 2 3 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 17 5 7 8 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
45 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 11 10 14 12 13 15 16 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 20 19 9 
3 1 2 18 
3 1 2 18 
31 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 13 15 14 12 16 
28 1 2 3 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 17 19 
7 1 2 3 20 9 18 9 
5 1 2 20 18 20 
30 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 14 15 12 13 16 
4 1 2 18 20 
47 1 2 3 9 9 9 9 9 4 9 9 6 5 7 8 9 10 5 17 7 8 10 10 10 10 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 22 16 12 15 13 14 16 
3 1 2 18 
30 1 2 3 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 14 13 12 15 16 
20 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 18 21 10 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
9 1 2 3 9 9 9 9 9 19 
7 1 2 3 20 9 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
19 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 19 17 10 
9 1 2 3 20 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 19 17 10 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 14 15 12 13 16 
33 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 19 17 10 
20 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 19 17 
4 1 2 18 20 
11 1 2 20 3 20 9 9 9 9 19 9 
20 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 14 15 13 12 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
22 1 2 3 20 9 9 4 5 6 7 8 9 10 10 11 10 16 14 15 12 13 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
25 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 14 15 12 13 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
5 1 2 3 19 9 
4 1 2 18 20 
3 1 2 18 
23 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 14 12 13 15 16 
6 1 2 3 9 18 9 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
9 1 2 3 9 9 9 9 18 9 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 10 11 10 15 14 12 13 16 
4 1 2 18 20 
5 1 2 23 18 23 
8 1 2 3 9 9 9 18 9 
3 1 2 18 
21 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 11 10 18 21 16 
4 1 2 18 20 
5 1 2 20 18 20 
17 1 2 3 4 5 6 7 8 9 11 10 16 14 15 13 12 16 
4 1 2 18 20 
5 1 2 3 19 9 
30 1 2 3 9 9 9 9 9 9 4 9 9 9 9 9 9 5 6 7 8 9 10 10 11 10 13 14 12 15 16 
5 1 2 23 18 23 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
19 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 18 21 16 
20 1 2 3 20 4 5 6 7 8 9 11 10 16 16 22 22 22 21 18 22 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
5 1 2 3 18 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
8 1 2 3 20 9 9 18 9 
20 1 2 3 9 9 9 4 6 5 7 8 9 11 10 16 15 12 14 13 16 
4 1 2 18 20 
5 1 2 20 18 20 
3 1 2 18 
20 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 20 18 20 
3 1 2 18 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
6 1 2 20 20 18 20 
5 1 2 3 19 9 
10 1 2 3 20 9 9 9 9 9 19 
22 1 2 3 20 9 4 6 5 7 8 9 10 10 10 11 10 16 14 13 12 15 16 
27 1 2 3 9 9 9 4 6 5 7 8 9 10 5 17 7 8 10 10 11 10 16 13 15 12 14 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
63 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 17 5 7 8 22 17 5 7 8 22 22 22 22 22 22 22 22 22 22 22 22 11 22 16 16 18 21 16 
28 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 14 13 15 12 16 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
28 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 17 5 7 8 16 14 15 13 12 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 19 9 
3 1 2 18 
5 1 2 23 18 23 
3 1 2 18 
5 1 2 20 18 20 
28 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 13 12 14 15 16 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 10 
6 1 2 20 20 18 20 
45 1 2 3 20 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 11 10 12 13 14 15 16 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
37 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 5 17 7 8 10 17 5 7 8 10 10 10 10 10 10 10 10 10 19 17 10 
11 1 2 3 20 9 9 9 9 9 9 19 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 15 13 12 16 
34 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
29 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 15 12 14 13 16 
35 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 14 13 12 15 16 
10 1 2 3 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
8 1 2 20 20 20 20 18 20 
5 1 2 20 18 20 
23 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
12 1 2 20 3 20 9 9 9 9 9 18 9 
5 1 2 20 18 20 
29 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
4 1 2 18 20 
20 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 13 14 15 12 16 
3 1 2 18 
3 1 2 18 
23 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
31 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
25 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 14 13 15 12 16 
4 1 2 18 20 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 17 19 
6 1 2 3 20 18 9 
8 1 2 20 20 3 20 19 9 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
5 1 2 20 18 20 
4 1 2 18 20 
5 1 2 20 18 20 
20 1 2 3 9 9 9 9 9 9 4 9 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
22 1 2 3 4 6 5 7 8 9 17 5 7 8 10 11 10 16 14 12 15 13 16 
3 1 2 18 
24 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 14 13 15 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 19 9 
17 1 2 3 9 4 6 5 7 8 9 10 10 11 10 18 21 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
7 1 2 20 3 20 18 9 
3 1 2 18 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
17 1 2 3 4 5 6 7 8 9 10 11 10 16 16 19 17 22 
26 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 17 19 10 
77 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 21 18 16 
3 1 2 18 
27 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 14 13 15 12 16 
4 1 2 18 20 
41 1 2 20 20 20 20 20 20 20 20 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 11 10 14 13 15 12 16 
4 1 2 18 20 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
6 1 2 20 20 18 20 
24 1 2 20 20 3 20 9 9 4 5 6 7 8 9 10 11 10 16 16 22 22 19 17 22 
5 1 2 20 18 20 
8 1 2 3 20 9 9 19 9 
4 1 2 18 20 
23 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 22 22 14 12 13 15 16 
33 1 2 20 20 3 20 9 9 9 4 6 5 7 8 9 10 11 10 5 17 7 8 16 22 22 22 11 22 14 12 13 15 16 
7 1 2 3 20 9 18 9 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
5 1 2 20 18 20 
21 1 2 20 3 20 9 4 5 6 7 8 9 11 10 16 16 14 12 15 13 16 
4 1 2 18 20 
12 1 2 3 20 9 9 9 9 9 9 18 9 
10 1 2 3 20 9 9 9 9 18 9 
5 1 2 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
27 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 14 12 13 15 16 
7 1 2 3 20 9 19 9 
4 1 2 18 20 
58 1 2 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 5 17 7 8 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
22 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
34 1 2 3 9 9 4 6 5 7 8 9 10 10 17 5 7 8 10 10 11 10 16 16 16 22 22 22 16 16 13 14 15 12 16 
21 1 2 3 20 9 4 5 6 7 8 9 10 10 10 11 10 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 20 9 4 5 6 7 8 9 11 10 21 18 16 
31 1 2 3 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
4 1 2 18 20 
24 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 11 10 16 16 14 13 15 12 16 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 21 18 16 
4 1 2 18 20 
8 1 2 3 20 9 9 19 9 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 15 13 12 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
25 1 2 20 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
24 1 2 3 9 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 10 10 10 19 17 
28 1 2 3 20 4 5 6 7 8 9 11 10 16 16 22 22 22 22 22 22 22 22 22 12 13 15 14 16 
3 1 2 18 
27 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 10 10 10 11 10 21 18 16 
16 1 2 3 4 5 6 7 8 9 11 10 14 13 15 12 16 
11 1 2 3 20 9 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
51 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 11 10 16 16 16 22 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 11 22 12 15 14 13 16 
3 1 2 18 
26 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 14 12 13 15 16 
27 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
34 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 16 16 22 22 13 14 12 15 16 
4 1 2 18 20 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 16 16 16 13 12 15 14 16 
6 1 2 23 23 18 23 
20 1 2 3 4 6 5 7 8 9 11 10 16 16 22 22 13 14 15 12 16 
18 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 18 21 10 
4 1 2 18 20 
3 1 2 18 
16 1 2 3 20 4 6 5 7 8 9 11 10 16 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
9 1 2 3 20 4 9 9 9 19 
3 1 2 18 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 10 10 11 10 21 18 16 
27 1 2 3 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 19 17 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
38 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 5 17 7 8 10 10 11 10 16 16 16 16 22 22 16 16 14 15 13 12 16 
7 1 2 3 9 9 19 9 
22 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 18 21 16 
3 1 2 18 
19 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 16 21 18 16 
22 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
52 1 2 3 20 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 17 5 7 8 10 10 10 10 10 17 5 7 8 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
19 1 2 3 9 4 6 5 7 8 9 10 11 10 16 14 12 13 15 16 
28 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
38 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 22 16 16 22 22 22 22 16 16 16 16 16 16 16 16 16 16 14 12 15 13 16 
26 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 16 16 14 13 12 15 16 
25 1 2 20 3 20 9 4 5 6 7 8 9 11 10 16 17 5 7 8 16 14 12 13 15 22 
36 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 14 12 15 13 16 
23 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 22 22 22 14 15 13 12 16 
3 1 2 18 
17 1 2 3 9 4 6 5 7 8 9 10 10 10 10 17 19 10 
24 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 11 10 12 14 13 15 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 12 13 15 16 
3 1 2 18 
5 1 2 20 18 20 
14 1 2 3 9 9 9 9 9 9 9 9 9 18 9 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
11 1 2 3 9 9 9 9 9 9 19 9 
6 1 2 3 4 19 9 
28 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 18 21 22 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
36 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 16 22 22 22 22 22 22 22 16 22 22 22 22 22 22 16 15 13 12 14 16 
3 1 2 18 
6 1 2 3 20 19 9 
18 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 18 21 16 
25 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 11 10 13 12 14 15 16 
19 1 2 3 9 4 5 6 7 8 9 10 11 10 16 14 12 13 15 16 
26 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 14 13 12 15 22 
3 1 2 18 
23 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 14 15 13 12 16 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 11 10 16 16 13 14 12 15 16 
3 1 2 18 
15 1 2 3 9 4 5 6 7 8 9 11 10 21 18 16 
30 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 16 22 22 18 21 22 
3 1 2 18 
5 1 2 3 19 9 
3 1 2 18 
29 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 11 10 16 16 14 13 15 12 16 
4 1 2 18 20 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 19 9 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 20 18 9 
5 1 2 3 18 9 
48 1 2 3 4 6 5 7 8 9 10 10 10 10 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 17 5 7 8 22 22 22 22 11 22 16 22 22 14 12 13 15 22 
6 1 2 3 20 19 9 
3 1 2 18 
5 1 2 20 18 20 
30 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
15 1 2 3 20 4 5 6 7 8 9 10 10 17 19 10 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
5 1 2 3 18 9 
7 1 2 3 9 9 18 9 
6 1 2 3 9 18 9 
28 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
7 1 2 3 20 9 18 9 
14 1 2 3 4 5 6 7 8 9 10 10 17 19 10 
20 1 2 3 4 5 6 7 8 9 11 10 16 16 22 16 15 13 12 14 16 
7 1 2 3 9 4 18 9 
4 1 2 18 20 
6 1 2 3 4 19 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
8 1 2 3 9 9 9 18 9 
22 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
7 1 2 3 4 9 19 9 
4 1 2 18 20 
7 1 2 20 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
8 1 2 20 3 20 9 18 9 
30 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 16 16 12 14 13 15 16 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
14 1 2 3 9 9 4 5 6 7 8 9 17 19 10 
30 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 5 17 7 8 10 10 11 10 12 13 15 14 16 
3 1 2 18 
32 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 11 10 16 18 21 16 
4 1 2 18 20 
4 1 2 18 20 
9 1 2 3 20 4 9 9 18 9 
14 1 2 3 20 4 6 5 7 8 9 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
21 1 2 3 20 9 9 4 5 6 7 8 9 10 5 17 7 8 10 18 21 10 
4 1 2 18 20 
3 1 2 18 
25 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 17 19 10 
21 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
38 1 2 3 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 10 10 11 10 16 5 17 7 8 16 14 13 15 12 22 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 22 18 21 22 
23 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 21 18 16 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
23 1 2 3 9 4 6 5 7 8 9 10 17 5 7 8 10 11 10 14 13 12 15 16 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 22 22 13 15 14 12 16 
6 1 2 3 20 18 9 
13 1 2 3 9 4 6 5 7 8 9 17 19 10 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
15 1 2 3 20 4 5 6 7 8 9 11 10 21 18 16 
3 1 2 18 
19 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 19 17 10 
27 1 2 3 20 9 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 22 22 14 13 12 15 16 
11 1 2 3 9 9 9 9 9 9 9 19 
18 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 17 19 10 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
30 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 22 22 13 14 15 12 16 
4 1 2 18 20 
23 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 11 10 13 14 12 15 16 
28 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 16 16 16 22 22 22 22 13 14 12 15 16 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 15 13 12 14 16 
14 1 2 3 9 9 9 9 9 9 9 9 9 19 9 
5 1 2 3 18 9 
16 1 2 3 4 6 5 7 8 9 11 10 14 15 13 12 16 
3 1 2 18 
7 1 2 3 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
29 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 13 14 12 15 16 
16 1 2 3 4 5 6 7 8 9 11 10 13 14 15 12 16 
4 1 2 18 20 
11 1 2 3 20 9 9 9 9 9 9 19 
4 1 2 18 20 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 14 12 15 13 16 
4 1 2 18 20 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
32 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 16 22 22 22 22 14 15 13 12 16 
43 1 2 3 20 9 4 6 5 7 8 9 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 14 15 13 12 16 
6 1 2 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 11 10 13 14 12 15 16 
35 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 5 17 7 8 10 10 11 10 16 18 21 16 
3 1 2 18 
24 1 2 3 9 9 9 9 4 5 6 7 8 9 11 10 16 22 22 22 13 12 14 15 16 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 14 13 12 15 16 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 17 19 10 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
7 1 2 3 20 4 18 9 
24 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 12 15 14 13 16 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 19 9 
28 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 5 17 7 8 16 12 15 13 14 22 
19 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 21 18 16 
16 1 2 3 9 9 9 9 4 6 5 7 8 9 18 21 10 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 20 18 20 
9 1 2 20 3 20 9 9 18 9 
8 1 2 3 20 9 9 18 9 
7 1 2 20 20 23 18 23 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 14 12 15 16 
26 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 16 16 22 22 22 14 13 15 12 16 
6 1 2 20 20 18 20 
6 1 2 3 9 19 9 
5 1 2 20 18 20 
18 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 4 19 9 
15 1 2 3 4 9 6 5 7 8 9 11 10 21 18 16 
29 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 15 13 12 14 16 
19 1 2 20 20 20 20 20 20 20 20 20 20 20 20 3 20 9 18 9 
11 1 2 20 20 3 20 9 9 9 18 9 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 15 12 13 16 
3 1 2 18 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 11 10 14 12 13 15 16 
4 1 2 18 20 
4 1 2 18 20 
10 1 2 3 9 9 9 9 9 9 19 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 19 17 10 
5 1 2 3 18 9 
4 1 2 18 20 
17 1 2 3 9 4 6 5 7 8 9 11 10 13 14 12 15 16 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 14 13 12 15 16 
29 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
8 1 2 3 9 9 9 19 9 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
10 1 2 3 9 9 9 9 9 9 19 
10 1 2 3 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 12 13 15 16 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 9 18 9 
3 1 2 18 
3 1 2 18 
40 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 5 17 7 8 16 14 13 15 12 22 
20 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 16 21 18 16 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
6 1 2 3 9 18 9 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
36 1 2 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 17 5 7 8 16 22 22 22 22 11 22 16 22 22 19 17 22 
3 1 2 18 
23 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 13 15 12 14 16 
5 1 2 20 18 20 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
3 1 2 18 
44 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 5 17 7 8 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
15 1 2 3 4 6 5 7 8 9 10 10 10 17 19 10 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
18 1 2 3 20 4 5 6 7 8 9 11 10 16 15 12 14 13 16 
3 1 2 18 
3 1 2 18 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
32 1 2 3 20 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 22 22 22 22 18 21 22 
17 1 2 3 9 9 4 5 6 7 8 9 10 11 10 18 21 16 
4 1 2 18 20 
3 1 2 18 
12 1 2 3 20 9 9 9 9 9 9 18 9 
35 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 11 10 16 16 22 22 22 22 19 17 22 
3 1 2 18 
9 1 2 3 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 4 9 18 9 
25 1 2 3 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 11 10 13 14 12 15 16 
4 1 2 18 20 
9 1 2 23 23 23 23 23 18 23 
3 1 2 18 
14 1 2 3 20 9 9 9 9 9 9 9 9 18 9 
60 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 17 5 7 8 16 22 22 22 22 22 22 22 22 11 22 16 16 14 13 12 15 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
58 1 2 3 20 9 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 16 16 17 5 7 8 16 14 13 12 15 22 
12 1 2 3 4 5 6 7 8 9 17 19 10 
34 1 2 3 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 11 10 18 21 16 
4 1 2 18 20 
22 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 11 10 16 22 19 17 22 
5 1 2 3 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
16 1 2 3 20 9 9 4 6 5 7 8 9 10 19 17 10 
7 1 2 3 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 14 12 13 15 22 
23 1 2 3 4 6 5 7 8 9 10 10 17 5 7 8 10 10 10 10 10 10 19 17 
3 1 2 18 
24 1 2 3 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 11 10 16 18 21 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
28 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 10 11 10 16 22 22 22 13 12 15 14 16 
4 1 2 18 20 
3 1 2 18 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 19 
33 1 2 3 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
22 1 2 3 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
34 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 22 19 17 22 
3 1 2 18 
40 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 16 22 22 22 22 22 22 16 16 16 16 16 22 22 22 22 22 22 22 14 15 13 12 16 
5 1 2 23 18 23 
3 1 2 18 
6 1 2 3 9 18 9 
5 1 2 20 18 20 
18 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 17 19 
18 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 17 19 10 
15 1 2 3 4 6 5 7 8 9 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
23 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 17 19 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
21 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 22 14 13 12 15 16 
36 1 2 3 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 22 17 5 7 8 22 22 22 11 22 14 12 13 15 16 
27 1 2 3 20 9 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 11 10 12 13 14 15 16 
31 1 2 3 9 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 22 16 22 22 22 16 21 18 16 
29 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 16 22 16 16 22 22 16 14 15 13 12 16 
4 1 2 18 20 
13 1 2 3 20 4 5 6 7 8 9 17 19 10 
48 1 2 3 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 17 5 7 8 10 10 11 10 16 22 22 22 22 22 22 14 12 13 15 16 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 17 5 7 8 10 11 10 12 13 14 15 16 
3 1 2 18 
4 1 2 18 20 
27 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 22 22 22 22 22 16 16 16 21 18 16 
16 1 2 3 4 5 6 7 8 9 10 10 11 10 21 18 16 
24 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 14 12 13 15 16 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
29 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 14 13 12 15 16 
3 1 2 18 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 11 10 18 21 16 
7 1 2 20 3 20 18 9 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
19 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
9 1 2 20 3 20 9 9 18 9 
3 1 2 18 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
5 1 2 3 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 14 12 15 16 
17 1 2 3 20 4 6 5 7 8 9 10 10 10 10 19 17 10 
6 1 2 3 9 19 9 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 18 9 
36 1 2 3 20 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 11 10 16 22 22 22 22 22 16 16 16 16 21 18 16 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 17 19 
3 1 2 18 
29 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 11 10 16 16 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
8 1 2 3 9 9 9 9 19 
3 1 2 18 
23 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
23 1 2 3 4 6 5 7 8 9 10 11 10 16 16 16 16 22 22 15 12 14 13 22 
3 1 2 18 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
27 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 9 9 9 19 
3 1 2 18 
34 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 16 22 22 22 22 22 22 14 12 15 13 16 
35 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 5 17 7 8 22 22 22 22 22 11 22 14 12 13 15 16 
4 1 2 18 20 
25 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
7 1 2 3 9 9 19 9 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
15 1 2 3 20 4 5 6 7 8 9 10 10 17 19 10 
4 1 2 18 20 
45 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 19 17 22 
15 1 2 3 4 6 5 7 8 9 10 10 10 19 17 10 
30 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 19 17 10 
40 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 14 13 12 15 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 13 12 15 16 
7 1 2 3 20 4 18 9 
6 1 2 3 20 19 9 
16 1 2 3 4 6 5 7 8 9 11 10 14 12 13 15 16 
28 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 12 14 13 15 16 
5 1 2 3 19 9 
4 1 2 18 20 
55 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 5 17 7 8 10 10 11 10 16 16 16 5 17 7 8 22 22 22 22 22 22 22 11 22 14 13 15 12 16 
3 1 2 18 
30 1 2 3 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 19 17 
7 1 2 3 20 9 18 9 
6 1 2 3 20 18 9 
16 1 2 3 4 5 6 7 8 9 11 10 14 13 12 15 16 
3 1 2 18 
17 1 2 3 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
33 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 16 16 16 16 22 22 22 22 15 14 12 13 16 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
16 1 2 3 9 4 6 5 7 8 9 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
6 1 2 3 4 19 9 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
22 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 22 22 14 15 13 12 22 
15 1 2 3 9 4 6 5 7 8 9 10 10 17 19 10 
5 1 2 3 18 9 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
17 1 2 3 9 9 9 4 5 6 7 8 9 10 10 18 21 10 
3 1 2 18 
9 1 2 20 20 20 3 20 19 9 
25 1 2 20 20 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 17 19 10 
6 1 2 3 20 19 9 
5 1 2 20 18 20 
3 1 2 18 
19 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
3 1 2 18 
6 1 2 3 9 19 9 
29 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 16 16 16 16 16 16 22 22 16 14 12 13 15 16 
3 1 2 18 
19 1 2 3 9 9 9 4 5 6 7 8 9 11 10 14 13 12 15 16 
54 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 17 5 7 8 10 10 11 10 16 16 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 12 14 13 15 16 
25 1 2 20 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 14 12 15 13 16 
34 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 21 18 16 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 21 18 16 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 11 10 18 21 16 
3 1 2 18 
10 1 2 3 9 9 9 9 9 19 9 
3 1 2 18 
15 1 2 3 4 6 5 7 8 9 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 18 9 
16 1 2 3 9 9 9 4 5 6 7 8 9 10 17 19 10 
20 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 17 19 10 
5 1 2 20 18 20 
47 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 16 16 22 22 22 22 22 17 5 7 8 16 22 22 22 22 22 5 17 7 8 22 22 22 22 22 15 14 12 13 22 
18 1 2 3 20 9 4 5 6 7 8 9 11 10 13 15 14 12 16 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
6 1 2 3 20 19 9 
4 1 2 18 20 
14 1 2 3 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
3 1 2 18 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 9 19 9 
4 1 2 18 20 
32 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 14 13 15 12 16 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 14 15 13 12 16 
4 1 2 18 20 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
4 1 2 18 20 
6 1 2 3 9 18 9 
4 1 2 18 20 
25 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 16 14 15 13 12 16 
27 1 2 3 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 13 12 14 15 16 
3 1 2 18 
5 1 2 3 18 9 
6 1 2 3 20 18 9 
3 1 2 18 
20 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 14 13 12 15 16 
5 1 2 20 18 20 
5 1 2 3 19 9 
4 1 2 18 20 
21 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
25 1 2 3 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 19 17 10 
5 1 2 3 19 9 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
32 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 16 22 22 22 22 22 22 14 15 13 12 16 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
14 1 2 3 4 5 6 7 8 9 10 10 17 19 10 
17 1 2 3 20 4 6 5 7 8 9 11 10 16 16 21 18 16 
27 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
17 1 2 3 20 4 5 6 7 8 9 11 10 14 13 12 15 16 
24 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 12 15 13 14 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
28 1 2 3 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 16 13 14 15 12 16 
3 1 2 18 
22 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 11 10 18 21 16 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
7 1 2 3 20 9 19 9 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 11 10 14 12 15 13 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 20 19 9 
42 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 16 16 13 14 12 15 16 
23 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 22 22 22 14 15 13 12 16 
4 1 2 18 20 
5 1 2 3 19 9 
7 1 2 20 3 20 18 9 
6 1 2 3 20 18 9 
6 1 2 3 20 18 9 
20 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
22 1 2 20 20 3 20 4 6 5 7 8 9 10 10 11 10 16 13 15 12 14 16 
32 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 22 22 22 16 16 22 22 22 22 22 22 22 13 14 15 12 16 
18 1 2 3 9 4 6 5 7 8 9 11 10 16 14 12 15 13 16 
5 1 2 20 18 20 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 9 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
25 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 22 22 14 13 15 12 16 
4 1 2 18 20 
17 1 2 20 3 20 4 6 5 7 8 9 10 10 10 17 19 10 
6 1 2 20 20 18 20 
3 1 2 18 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
13 1 2 3 20 9 9 9 9 9 9 9 19 9 
16 1 2 3 20 4 5 6 7 8 9 10 10 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
28 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 18 21 16 
4 1 2 18 20 
22 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 16 21 18 16 
4 1 2 18 20 
23 1 2 20 20 3 20 4 6 5 7 8 9 10 10 10 10 11 10 12 14 13 15 16 
31 1 2 3 20 9 9 9 4 6 5 7 8 9 11 10 16 16 16 16 16 16 16 16 16 16 16 13 14 12 15 16 
27 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 11 10 13 15 12 14 16 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
42 1 2 3 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 16 22 22 22 22 22 22 22 22 15 13 14 12 16 
4 1 2 18 20 
23 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 21 18 16 
5 1 2 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
6 1 2 20 20 18 20 
5 1 2 3 19 9 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
49 1 2 3 9 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 10 10 17 5 7 8 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 16 12 13 15 14 16 
18 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 19 17 
25 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 16 16 16 16 16 16 18 21 16 
18 1 2 3 9 4 9 6 5 7 8 9 10 11 10 16 21 18 16 
5 1 2 20 18 20 
12 1 2 3 4 5 6 7 8 9 19 17 10 
14 1 2 3 4 6 5 7 8 9 11 10 18 21 16 
6 1 2 3 20 18 9 
4 1 2 18 20 
18 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 19 17 10 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
28 1 2 3 4 5 6 7 8 9 5 17 7 8 10 11 10 16 16 22 22 22 22 22 14 13 15 12 16 
28 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 22 18 21 22 
4 1 2 18 20 
16 1 2 3 4 5 6 7 8 9 11 10 14 15 13 12 16 
4 1 2 18 20 
54 1 2 3 20 4 5 6 7 8 9 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 13 14 15 12 16 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 17 19 10 
6 1 2 20 20 18 20 
20 1 2 3 4 6 5 7 8 9 11 10 16 16 22 16 14 13 12 15 16 
11 1 2 3 9 9 9 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
38 1 2 3 20 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 11 10 16 16 16 16 16 16 16 16 17 19 16 
3 1 2 18 
6 1 2 3 20 18 9 
29 1 2 3 9 9 4 6 5 7 8 9 10 10 10 5 17 7 8 10 10 10 10 11 10 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
5 1 2 3 19 9 
5 1 2 3 18 9 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
30 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 16 16 22 22 22 22 13 14 12 15 16 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
31 1 2 3 20 9 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 11 10 16 16 22 22 22 21 18 16 
7 1 2 3 20 9 18 9 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
3 1 2 18 
6 1 2 3 20 19 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 18 9 
21 1 2 3 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 19 17 10 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
41 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 11 10 14 15 13 12 16 
16 1 2 3 9 4 6 5 7 8 9 10 10 10 10 19 17 
30 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 16 22 22 22 16 22 22 22 22 14 12 13 15 16 
5 1 2 3 18 9 
15 1 2 3 9 4 5 6 7 8 9 10 10 17 19 10 
4 1 2 18 20 
21 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 17 19 10 
28 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
21 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
7 1 2 20 3 20 18 9 
4 1 2 18 20 
46 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 17 5 7 8 22 22 22 22 11 22 16 22 22 22 22 22 22 14 13 15 12 16 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
23 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 16 14 12 13 15 16 
14 1 2 3 9 9 9 9 9 9 9 9 9 19 9 
6 1 2 3 20 18 9 
35 1 2 3 20 9 9 9 4 6 5 7 8 9 11 10 16 16 16 22 22 16 22 22 22 22 22 22 22 22 16 15 13 12 14 16 
3 1 2 18 
33 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 21 18 16 
4 1 2 18 20 
6 1 2 3 20 19 9 
35 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 22 22 22 22 22 22 22 16 16 13 14 15 12 16 
4 1 2 18 20 
10 1 2 3 9 9 9 9 9 9 19 
6 1 2 3 9 18 9 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
23 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
4 1 2 18 20 
27 1 2 3 20 9 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 16 13 14 15 12 16 
56 1 2 20 3 20 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 16 16 16 22 16 22 22 22 17 5 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
20 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 11 10 16 22 22 16 14 12 13 15 16 
4 1 2 18 20 
20 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 17 19 
23 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 21 18 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
24 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
17 1 2 3 9 4 5 6 7 8 9 10 11 10 16 18 21 22 
3 1 2 18 
35 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 21 18 16 
4 1 2 18 20 
30 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 11 10 18 21 16 
26 1 2 3 20 9 9 4 5 6 7 8 9 10 10 11 10 16 16 16 22 22 12 14 13 15 16 
4 1 2 18 20 
5 1 2 3 18 9 
48 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 12 14 13 15 16 
22 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 22 22 15 13 12 14 16 
3 1 2 18 
4 1 2 18 20 
27 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 11 10 13 14 12 15 16 
33 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 21 18 16 
22 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 16 22 22 16 18 21 16 
6 1 2 20 20 18 20 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
16 1 2 3 4 5 6 7 8 9 10 11 10 16 18 21 16 
21 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 16 14 12 13 15 16 
40 1 2 3 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 14 13 15 12 16 
3 1 2 18 
40 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
11 1 2 3 20 9 9 9 9 9 18 9 
43 1 2 3 9 9 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 5 17 7 8 10 10 10 5 17 7 8 10 10 10 10 10 10 19 17 
5 1 2 20 18 20 
7 1 2 23 23 23 18 23 
23 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 16 22 22 14 13 15 12 16 
31 1 2 3 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 11 10 16 22 16 16 13 15 14 12 16 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 14 13 12 15 16 
23 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 18 21 16 
3 1 2 18 
25 1 2 3 9 4 6 5 7 8 9 10 10 10 10 17 5 7 8 10 10 11 10 21 18 16 
6 1 2 20 20 18 20 
4 1 2 18 20 
29 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 18 21 16 
16 1 2 3 20 4 6 5 7 8 9 10 10 10 17 19 10 
3 1 2 18 
29 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 18 21 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 14 13 15 12 16 
29 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 21 18 16 
18 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 19 17 10 
9 1 2 3 20 9 9 9 9 19 
9 1 2 3 20 9 9 9 18 9 
60 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 17 19 16 
6 1 2 20 20 18 20 
16 1 2 3 20 9 4 6 5 7 8 9 10 10 10 17 19 
18 1 2 3 20 4 6 5 7 8 9 10 11 10 13 14 12 15 16 
3 1 2 18 
32 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 17 19 10 
10 1 2 3 20 9 9 9 9 18 9 
24 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 10 11 10 14 12 13 15 16 
23 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 18 21 16 
28 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 11 10 13 14 12 15 16 
5 1 2 3 18 9 
30 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 5 17 7 8 10 10 11 10 14 13 12 15 16 
7 1 2 3 9 9 9 19 
10 1 2 20 20 3 20 9 9 18 9 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 15 12 13 14 16 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 22 14 13 12 15 16 
3 1 2 18 
32 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
9 1 2 3 9 9 9 9 19 9 
25 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 14 13 15 12 16 
4 1 2 18 20 
3 1 2 18 
40 1 2 3 4 6 5 7 8 9 17 5 7 8 10 17 5 7 8 10 10 10 10 10 10 10 10 11 10 16 22 22 22 16 16 16 14 13 15 12 16 
6 1 2 3 9 18 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
34 1 2 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 11 10 16 22 22 16 22 22 22 16 14 13 12 15 16 
3 1 2 18 
25 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 13 14 12 15 16 
5 1 2 20 18 20 
20 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 13 14 12 15 16 
6 1 2 3 20 19 9 
37 1 2 20 3 20 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 17 5 7 8 16 22 22 22 22 22 11 22 13 14 15 12 16 
6 1 2 3 20 19 9 
32 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 11 10 16 16 16 22 16 22 19 17 22 
35 1 2 3 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 16 22 22 22 22 22 22 22 22 22 16 21 18 16 
21 1 2 3 4 6 5 7 8 9 5 17 7 8 10 11 10 14 12 13 15 16 
3 1 2 18 
9 1 2 3 9 4 9 9 9 19 
45 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 16 16 16 16 22 22 22 22 17 5 7 8 22 22 22 22 11 22 16 16 16 22 12 13 14 15 16 
21 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 18 21 16 
15 1 2 3 4 6 5 7 8 9 10 10 10 17 19 10 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
22 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 14 12 13 15 16 
6 1 2 3 20 18 9 
3 1 2 18 
6 1 2 3 9 19 9 
5 1 2 20 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
27 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 16 22 22 22 21 18 16 
21 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
14 1 2 3 4 5 6 7 8 9 10 10 17 19 10 
33 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 19 17 10 
3 1 2 18 
29 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 11 10 5 17 7 8 16 22 14 12 13 15 22 
34 1 2 3 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
4 1 2 18 20 
8 1 2 3 9 9 9 19 9 
3 1 2 18 
55 1 2 3 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 17 5 7 8 10 17 5 7 8 10 10 10 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 14 12 13 15 16 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
27 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 16 16 22 22 22 22 22 12 13 14 15 16 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 16 22 21 18 22 
3 1 2 18 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 13 14 15 12 16 
16 1 2 3 9 9 9 4 6 5 7 8 9 10 19 17 10 
28 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 17 5 7 8 10 10 10 11 10 18 21 16 
52 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 16 22 16 16 16 21 18 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
9 1 2 3 20 9 9 9 18 9 
4 1 2 18 20 
5 1 2 3 18 9 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 14 13 15 12 16 
5 1 2 3 18 9 
11 1 2 3 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 4 18 9 
9 1 2 3 20 9 9 9 18 9 
39 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 17 5 7 8 10 17 5 7 8 10 10 10 10 10 11 10 13 14 15 12 16 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 10 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
20 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 16 18 21 16 
36 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
8 1 2 20 3 20 9 18 9 
40 1 2 3 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 16 16 16 22 22 22 22 22 22 22 22 22 16 13 14 12 15 16 
3 1 2 18 
4 1 2 18 20 
9 1 2 3 20 9 9 9 9 19 
3 1 2 18 
5 1 2 20 18 20 
21 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 13 14 15 12 16 
3 1 2 18 
40 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 19 17 22 
25 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
5 1 2 3 9 19 
3 1 2 18 
3 1 2 18 
23 1 2 20 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 17 19 10 
67 1 2 3 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 12 13 15 14 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
25 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 16 13 14 15 12 16 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 12 13 15 16 
13 1 2 3 9 4 6 5 7 8 9 17 19 10 
71 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 17 19 
3 1 2 18 
23 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 16 16 16 14 13 15 12 16 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 19 9 
10 1 2 3 20 9 9 9 9 9 19 
6 1 2 3 9 19 9 
3 1 2 18 
25 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
18 1 2 3 20 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
4 1 2 18 20 
7 1 2 3 9 9 19 9 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
4 1 2 18 20 
24 1 2 3 20 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 18 21 16 
3 1 2 18 
4 1 2 18 20 
5 1 2 3 18 9 
8 1 2 20 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
31 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 17 5 7 8 10 10 10 10 10 11 10 14 12 13 15 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
28 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 14 12 13 15 16 
26 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 16 14 13 15 12 16 
21 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 10 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
3 1 2 18 
5 1 2 20 18 20 
28 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 16 22 22 22 22 22 22 16 13 14 12 15 16 
26 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
5 1 2 3 19 9 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
45 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 17 5 7 8 10 10 10 11 10 16 22 17 5 7 8 22 22 22 22 22 22 22 22 11 22 14 12 13 15 16 
19 1 2 3 9 4 6 5 7 8 9 10 11 10 16 14 13 15 12 16 
16 1 2 3 20 9 4 5 6 7 8 9 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
17 1 2 3 9 9 4 6 5 7 8 9 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 20 18 9 
12 1 2 3 4 6 5 7 8 9 10 17 19 
22 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 10 
17 1 2 3 4 5 6 7 8 9 11 10 16 22 22 21 18 22 
6 1 2 3 9 19 9 
3 1 2 18 
26 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 17 5 7 8 16 13 12 14 15 22 
29 1 2 3 20 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
6 1 2 20 20 18 20 
22 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 14 15 13 12 16 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 13 12 14 15 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 14 12 15 16 
17 1 2 3 4 5 6 7 8 9 11 10 16 13 12 14 15 16 
3 1 2 18 
32 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
37 1 2 3 20 4 5 6 7 8 9 10 10 10 10 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 16 16 16 14 12 13 15 16 
32 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 16 16 16 22 22 14 13 12 15 22 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
44 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 11 10 16 22 22 22 5 17 7 8 16 12 14 13 15 22 
39 1 2 3 9 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 16 21 18 22 
4 1 2 18 20 
3 1 2 18 
30 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 11 10 16 22 22 22 22 22 13 12 14 15 16 
6 1 2 3 20 18 9 
3 1 2 18 
32 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 5 17 7 8 10 10 11 10 16 16 16 22 22 21 18 22 
12 1 2 3 4 5 6 7 8 9 19 17 10 
23 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 22 18 21 16 
3 1 2 18 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
31 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 22 22 14 12 13 15 16 
25 1 2 3 9 9 9 4 6 5 7 8 9 10 10 17 5 7 8 10 10 11 10 18 21 16 
22 1 2 3 20 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
27 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 17 19 10 
42 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 17 5 7 8 10 17 5 7 8 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
9 1 2 3 9 9 9 9 19 9 
3 1 2 18 
5 1 2 3 18 9 
5 1 2 3 18 9 
66 1 2 3 9 9 9 4 9 9 9 5 6 7 8 9 10 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 22 22 16 22 22 22 22 22 14 15 13 12 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 11 10 21 18 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
37 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 16 16 17 5 7 8 16 13 14 15 12 22 
31 1 2 3 9 9 9 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
24 1 2 3 20 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 10 17 19 10 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 18 21 16 
24 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 11 10 21 18 16 
5 1 2 3 19 9 
19 1 2 3 20 4 5 6 7 8 9 10 11 10 16 14 12 13 15 16 
39 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 16 22 22 16 16 22 22 22 22 16 5 17 7 8 16 14 13 15 12 22 
28 1 2 20 3 20 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 16 16 16 16 21 18 16 
20 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 16 21 18 16 
3 1 2 18 
24 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 19 17 10 
4 1 2 18 20 
29 1 2 3 20 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 16 16 13 12 14 15 16 
7 1 2 3 20 9 18 9 
3 1 2 18 
9 1 2 3 20 9 9 9 19 9 
22 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 22 22 14 13 12 15 16 
3 1 2 18 
22 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
35 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
7 1 2 23 23 23 18 23 
58 1 2 3 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 15 13 12 14 16 
55 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 5 17 7 8 10 10 5 17 7 8 10 10 5 17 7 8 10 10 17 5 7 8 10 10 10 10 11 10 16 16 16 16 16 16 16 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
7 1 2 3 20 9 18 9 
19 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 19 17 10 
19 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 22 19 17 22 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
82 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 17 19 22 
7 1 2 3 20 9 18 9 
5 1 2 3 18 9 
15 1 2 3 9 4 5 6 7 8 9 10 10 17 19 10 
21 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 19 17 10 
23 1 2 3 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 14 12 13 15 16 
3 1 2 18 
6 1 2 3 20 18 9 
37 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 22 16 16 5 17 7 8 16 14 12 13 15 22 
6 1 2 3 9 18 9 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
23 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 11 10 12 15 14 13 16 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 15 12 13 14 16 
3 1 2 18 
11 1 2 20 3 20 9 9 9 9 9 19 
15 1 2 3 20 4 6 5 7 8 9 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
29 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 16 16 22 22 14 13 15 12 16 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 20 9 4 6 5 7 8 9 10 10 10 11 10 14 13 15 12 16 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 17 19 10 
23 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
6 1 2 3 9 19 9 
5 1 2 20 18 20 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 18 9 
4 1 2 18 20 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 18 9 
4 1 2 18 20 
22 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 14 13 15 12 16 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 11 10 21 18 16 
9 1 2 3 20 9 9 9 18 9 
4 1 2 18 20 
28 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 22 22 22 16 15 14 12 13 16 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
9 1 2 3 9 9 9 9 18 9 
5 1 2 3 18 9 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
34 1 2 20 3 20 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 22 22 22 22 5 17 7 8 16 15 13 12 14 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
23 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 18 21 16 
3 1 2 18 
19 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
5 1 2 23 18 23 
21 1 2 3 4 9 5 6 7 8 9 10 10 10 11 10 16 14 13 15 12 16 
3 1 2 18 
22 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
5 1 2 23 18 23 
3 1 2 18 
44 1 2 3 20 9 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 17 5 7 8 10 10 10 10 10 10 10 11 10 16 16 16 22 22 22 14 12 13 15 16 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
19 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 17 19 10 
13 1 2 3 20 9 9 9 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
14 1 2 3 20 9 4 5 6 7 8 9 19 17 10 
26 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
11 1 2 3 9 9 9 9 9 9 19 9 
39 1 2 20 3 20 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
3 1 2 18 
14 1 2 3 20 9 4 6 5 7 8 9 19 17 10 
3 1 2 18 
3 1 2 18 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 5 17 7 8 10 11 10 14 12 15 13 16 
58 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 22 22 22 22 22 22 22 11 22 5 17 7 8 16 14 12 15 13 22 
29 1 2 20 3 20 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 11 10 16 16 22 22 18 21 16 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 3 19 9 
3 1 2 18 
6 1 2 3 9 19 9 
31 1 2 3 20 9 4 5 6 7 8 9 10 10 17 5 7 8 10 11 10 16 16 22 22 16 16 14 12 13 15 16 
3 1 2 18 
5 1 2 20 18 20 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 19 17 16 
3 1 2 18 
7 1 2 3 9 9 19 9 
40 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 11 10 17 5 7 8 16 22 22 22 22 22 22 22 22 22 11 22 14 13 15 12 16 
3 1 2 18 
40 1 2 3 20 9 9 4 9 6 5 7 8 9 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 11 10 16 22 22 22 22 21 18 22 
3 1 2 18 
39 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 16 16 21 18 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 19 17 10 
32 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 16 16 22 22 22 16 22 17 19 22 
3 1 2 18 
6 1 2 3 9 18 9 
33 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 11 10 16 22 22 22 18 21 16 
5 1 2 3 18 9 
9 1 2 3 20 9 9 9 9 19 
19 1 2 3 9 9 4 5 6 7 8 9 10 11 10 14 15 13 12 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 19 9 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 19 9 
27 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 15 14 12 13 22 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
17 1 2 3 4 5 6 7 8 9 11 10 16 14 15 13 12 16 
6 1 2 3 9 18 9 
5 1 2 3 18 9 
5 1 2 3 18 9 
38 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 17 19 
17 1 2 3 9 9 4 5 6 7 8 9 11 10 16 18 21 16 
19 1 2 3 4 6 5 7 8 9 10 10 10 11 10 14 12 13 15 16 
5 1 2 23 18 23 
7 1 2 3 20 9 18 9 
3 1 2 18 
19 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 21 18 16 
7 1 2 3 20 9 19 9 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 13 14 12 15 16 
11 1 2 3 9 9 9 9 9 9 19 9 
5 1 2 3 18 9 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 11 10 16 22 16 18 21 16 
24 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 17 19 10 
12 1 2 3 4 5 6 7 8 9 19 17 10 
3 1 2 18 
3 1 2 18 
25 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 9 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 17 19 
13 1 2 3 20 4 5 6 7 8 9 18 21 10 
4 1 2 18 20 
4 1 2 18 20 
29 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 16 16 21 18 16 
7 1 2 20 3 20 18 9 
21 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 19 
27 1 2 3 9 4 5 6 7 8 9 10 11 10 5 17 7 8 16 22 22 22 22 22 22 21 18 22 
17 1 2 3 20 4 6 5 7 8 9 11 10 13 12 15 14 16 
4 1 2 18 20 
25 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 15 13 12 16 
3 1 2 18 
5 1 2 3 18 9 
27 1 2 3 9 4 5 6 7 8 9 11 10 16 16 16 22 22 22 22 16 22 22 14 12 13 15 16 
5 1 2 3 19 9 
5 1 2 3 18 9 
28 1 2 20 3 20 9 9 4 6 5 7 8 9 10 11 10 16 22 22 16 22 22 16 14 13 12 15 16 
3 1 2 18 
6 1 2 3 9 18 9 
22 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 17 19 
31 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 5 17 7 8 16 12 13 14 15 22 
3 1 2 18 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 19 17 10 
6 1 2 3 9 18 9 
6 1 2 3 20 18 9 
3 1 2 18 
6 1 2 23 23 18 23 
4 1 2 18 20 
25 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 11 10 16 16 21 18 16 
4 1 2 18 20 
5 1 2 3 18 9 
37 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
8 1 2 3 9 9 9 19 9 
15 1 2 3 9 9 4 6 5 7 8 9 10 19 17 10 
6 1 2 3 20 18 9 
4 1 2 18 20 
32 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 16 16 18 21 16 
21 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
30 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 16 16 16 16 16 22 14 12 13 15 16 
3 1 2 18 
27 1 2 3 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 11 10 18 21 16 
4 1 2 18 20 
28 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 13 14 15 12 22 
21 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 17 19 10 
27 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 16 14 12 13 15 16 
5 1 2 3 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
16 1 2 3 9 9 4 6 5 7 8 9 10 10 19 17 10 
3 1 2 18 
7 1 2 3 9 9 19 9 
23 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 10 
16 1 2 3 20 9 4 6 5 7 8 9 10 10 17 19 10 
9 1 2 3 9 9 9 9 19 9 
9 1 2 3 9 9 9 9 19 9 
31 1 2 20 20 3 20 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 10 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 17 19 10 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 13 14 15 12 16 
29 1 2 3 4 6 5 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 16 22 22 14 13 12 15 16 
3 1 2 18 
17 1 2 3 20 4 5 6 7 8 9 10 10 10 10 17 19 10 
22 1 2 20 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 18 21 10 
22 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 16 14 12 13 15 16 
4 1 2 18 20 
4 1 2 18 20 
9 1 2 3 20 9 9 9 18 9 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 14 12 13 15 16 
3 1 2 18 
24 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 14 12 13 15 16 
44 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 16 22 22 22 22 16 17 5 7 8 22 22 22 22 22 22 22 22 11 22 15 14 12 13 16 
32 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 11 10 17 5 7 8 16 14 15 13 12 22 
3 1 2 18 
8 1 2 3 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
21 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 15 13 14 12 22 
32 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 19 17 
29 1 2 20 3 20 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
38 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 16 22 14 12 13 15 22 
3 1 2 18 
7 1 2 3 9 9 19 9 
11 1 2 3 9 9 9 9 9 9 18 9 
13 1 2 3 9 9 9 9 9 9 9 9 18 9 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
52 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 16 16 16 16 16 22 22 22 22 22 22 22 22 22 16 16 5 17 7 8 16 13 14 12 15 22 
12 1 2 3 9 9 9 9 9 9 9 19 9 
3 1 2 18 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 17 5 7 8 10 10 10 19 17 10 
3 1 2 18 
43 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 16 16 22 22 22 16 16 22 5 17 7 8 22 22 22 22 22 22 22 17 19 22 
3 1 2 18 
33 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 11 10 16 16 16 22 22 22 22 22 21 18 16 
23 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 14 12 15 13 16 
4 1 2 18 20 
24 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
49 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 22 22 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 16 12 13 14 15 16 
3 1 2 18 
28 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 9 19 9 
3 1 2 18 
17 1 2 3 20 9 4 6 5 7 8 9 10 10 10 19 17 10 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 13 12 15 16 
29 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
19 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 17 19 10 
28 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 12 13 15 14 16 
48 1 2 3 20 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 17 5 7 8 10 10 10 10 11 10 16 14 12 15 13 16 
28 1 2 3 4 5 6 7 8 9 10 10 11 10 16 23 16 22 22 22 22 22 22 22 14 15 13 12 16 
3 1 2 18 
3 1 2 18 
25 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 10 17 
33 1 2 3 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
25 1 2 3 20 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 11 10 21 18 16 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
22 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 11 10 14 12 13 15 16 
22 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 13 14 15 12 16 
3 1 2 18 
28 1 2 3 4 9 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
3 1 2 18 
28 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 11 10 16 16 12 14 13 15 16 
3 1 2 18 
14 1 2 3 9 9 4 5 6 7 8 9 17 19 10 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
15 1 2 3 20 9 4 5 6 7 8 9 10 19 17 10 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
3 1 2 18 
5 1 2 20 18 20 
24 1 2 3 9 9 9 4 6 5 7 8 9 11 10 16 22 22 22 22 14 13 15 12 22 
21 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 17 19 10 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
28 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 5 17 7 8 10 10 10 11 10 21 18 16 
4 1 2 18 20 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
6 1 2 3 20 19 9 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
25 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 17 5 7 8 10 18 21 10 
4 1 2 18 20 
6 1 2 3 9 19 9 
5 1 2 3 19 9 
6 1 2 3 9 19 9 
32 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 11 10 16 16 16 22 19 17 22 
3 1 2 18 
5 1 2 3 19 9 
8 1 2 3 20 9 9 18 9 
7 1 2 3 9 9 18 9 
4 1 2 18 20 
8 1 2 3 20 9 9 9 19 
3 1 2 18 
4 1 2 18 20 
5 1 2 3 19 9 
7 1 2 3 9 9 18 9 
3 1 2 18 
32 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
8 1 2 3 9 9 9 19 9 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
16 1 2 3 4 5 6 7 8 9 11 10 14 13 15 12 16 
18 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 21 18 16 
18 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 19 17 10 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
22 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 18 21 16 
18 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 21 18 16 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 10 10 11 10 14 13 12 15 16 
20 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 14 15 13 12 16 
4 1 2 18 20 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 16 18 21 16 
24 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 16 14 12 13 15 16 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
3 1 2 18 
21 1 2 3 20 9 4 5 6 7 8 9 10 5 17 7 8 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 14 15 13 12 16 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
21 1 2 20 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 19 17 10 
5 1 2 20 18 20 
4 1 2 18 20 
10 1 2 20 3 20 9 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
41 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
42 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 11 10 16 22 5 17 7 8 22 22 22 22 22 22 11 22 14 15 13 12 16 
5 1 2 3 19 9 
5 1 2 3 18 9 
24 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 10 17 
19 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 16 21 18 16 
3 1 2 18 
7 1 2 3 9 9 19 9 
24 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 15 13 14 12 16 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
16 1 2 3 20 9 4 6 5 7 8 9 10 10 19 17 10 
11 1 2 3 9 9 9 9 9 9 19 9 
23 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 13 14 15 12 16 
7 1 2 3 9 9 18 9 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 13 15 12 16 
13 1 2 3 20 9 9 9 9 9 9 9 19 9 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 19 17 
6 1 2 3 9 19 9 
5 1 2 20 18 20 
6 1 2 3 4 19 9 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 19 9 
15 1 2 3 4 5 6 7 8 9 10 11 10 21 18 16 
17 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 18 9 
5 1 2 3 18 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
25 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 21 18 16 
3 1 2 18 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
19 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 19 17 
28 1 2 3 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
23 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 15 14 12 13 16 
5 1 2 3 19 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
31 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 11 10 16 16 22 22 22 14 12 13 15 16 
19 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
20 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 19 17 
4 1 2 18 20 
5 1 2 3 19 9 
5 1 2 3 18 9 
7 1 2 3 9 9 19 9 
6 1 2 3 9 19 9 
3 1 2 18 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 21 18 16 
22 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 16 14 15 13 12 16 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 10 
38 1 2 3 20 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
21 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 19 17 10 
3 1 2 18 
7 1 2 3 20 9 18 9 
23 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 13 15 14 12 16 
6 1 2 3 9 18 9 
12 1 2 3 20 9 9 9 9 9 9 9 19 
26 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 13 14 12 15 16 
28 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 17 5 7 8 10 10 10 10 17 19 10 
6 1 2 3 9 19 9 
3 1 2 18 
22 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 10 11 10 21 18 16 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 15 13 12 14 16 
3 1 2 18 
4 1 2 18 20 
28 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 22 13 14 12 15 22 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
30 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 19 9 
25 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
5 1 2 20 18 20 
3 1 2 18 
14 1 2 20 3 20 9 9 9 9 9 9 9 9 19 
7 1 2 3 20 9 19 9 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 19 17 
4 1 2 18 20 
22 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
19 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
3 1 2 18 
14 1 2 3 20 9 9 9 9 9 9 9 9 18 9 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 21 18 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 15 13 14 12 16 
3 1 2 18 
26 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 16 13 14 15 12 16 
4 1 2 18 20 
7 1 2 20 3 20 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
25 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 14 13 15 12 16 
4 1 2 18 20 
22 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
22 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 14 12 13 15 16 
11 1 2 3 9 9 9 9 9 9 9 19 
5 1 2 3 18 9 
5 1 2 3 18 9 
22 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 11 10 14 13 15 12 16 
13 1 2 3 20 9 9 9 9 9 9 9 9 19 
28 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 21 18 16 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 15 13 12 16 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
7 1 2 20 20 20 20 19 
31 1 2 3 9 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 11 10 16 22 22 22 22 15 14 12 13 16 
3 1 2 18 
19 1 2 3 9 4 6 5 7 8 9 10 10 11 10 13 12 14 15 16 
4 1 2 18 20 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
19 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
6 1 2 3 9 19 9 
4 1 2 18 20 
31 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 16 16 16 22 22 22 22 12 14 13 15 16 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
24 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 16 12 14 13 15 16 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 18 9 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
27 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 16 16 22 12 14 13 15 16 
32 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
21 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
30 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 13 14 15 12 16 
31 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 16 17 5 7 8 16 22 22 22 11 22 13 14 15 12 16 
23 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 14 15 13 12 16 
23 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
27 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 16 14 15 13 12 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 12 15 13 14 16 
4 1 2 18 20 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
25 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 16 12 13 14 15 16 
4 1 2 18 20 
3 1 2 18 
26 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 22 19 17 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 17 19 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
19 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 19 17 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
29 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 19 17 
11 1 2 3 20 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
16 1 2 3 9 4 6 5 7 8 9 10 11 10 21 18 16 
4 1 2 18 20 
4 1 2 18 20 
7 1 2 3 20 9 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
18 1 2 3 20 9 4 6 5 7 8 9 11 10 14 13 12 15 16 
4 1 2 18 20 
3 1 2 18 
24 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
9 1 2 3 20 9 9 9 19 9 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
13 1 2 3 20 4 5 6 7 8 9 17 19 10 
3 1 2 18 
6 1 2 3 9 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
45 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 14 12 13 15 16 
5 1 2 3 19 9 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
27 1 2 20 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 19 17 10 
6 1 2 3 9 19 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
6 1 2 3 20 18 9 
37 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 22 22 14 13 12 15 16 
4 1 2 18 20 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
31 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 16 16 16 22 22 22 18 21 16 
8 1 2 3 20 9 9 18 9 
25 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
6 1 2 3 9 19 9 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 9 19 
24 1 2 3 9 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 14 15 13 12 16 
19 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
4 1 2 18 20 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 19 17 
25 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 11 10 13 14 12 15 16 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 13 15 14 12 16 
3 1 2 18 
5 1 2 20 18 20 
4 1 2 18 20 
7 1 2 3 9 9 18 9 
4 1 2 18 20 
42 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 17 5 7 8 22 22 22 22 22 22 22 22 22 22 11 22 16 22 16 13 14 12 15 16 
4 1 2 18 20 
34 1 2 3 4 6 5 7 8 9 10 10 10 17 5 7 8 10 11 10 16 22 22 16 16 22 22 22 22 22 14 12 15 13 16 
3 1 2 18 
43 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 16 16 17 5 7 8 16 13 14 12 15 22 
14 1 2 3 20 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
7 1 2 3 9 9 18 9 
3 1 2 18 
6 1 2 20 20 18 20 
12 1 2 3 4 5 6 7 8 9 21 18 10 
11 1 2 3 20 9 9 9 9 9 18 9 
24 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
5 1 2 3 18 9 
28 1 2 3 9 9 4 5 6 7 8 9 11 10 17 5 7 8 16 22 22 22 11 22 15 13 12 14 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
66 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 5 17 7 8 10 10 11 10 5 17 7 8 16 11 22 16 22 22 22 22 22 22 22 22 22 22 16 16 22 5 17 7 8 22 22 22 22 22 22 22 22 22 11 22 16 13 12 14 15 16 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
19 1 2 3 9 4 6 5 7 8 9 10 10 11 10 14 12 15 13 16 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
8 1 2 3 20 9 9 18 9 
16 1 2 3 20 4 6 5 7 8 9 10 10 10 10 17 19 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 17 19 10 
23 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 13 12 14 15 16 
21 1 2 3 20 9 4 5 6 7 8 9 10 10 10 11 10 15 13 12 14 16 
37 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 13 14 12 15 16 
14 1 2 3 9 9 4 6 5 7 8 9 17 19 10 
29 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 5 17 7 8 10 10 11 10 16 18 21 16 
8 1 2 20 20 3 20 18 9 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 11 10 16 18 21 16 
9 1 2 3 20 9 9 9 19 9 
5 1 2 3 19 9 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 15 13 12 14 16 
17 1 2 3 4 5 6 7 8 9 10 11 10 15 14 12 13 16 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 4 9 19 9 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 19 9 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 13 15 12 16 
7 1 2 3 20 9 18 9 
24 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
25 1 2 23 23 20 23 23 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
7 1 2 3 20 9 18 9 
25 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
27 1 2 23 23 20 23 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
7 1 2 3 20 9 18 9 
3 1 2 18 
19 1 2 3 9 4 5 6 7 8 9 11 10 16 16 14 15 13 12 16 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 14 15 13 12 16 
40 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 11 10 18 21 16 
20 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 13 15 12 14 16 
40 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 16 21 18 16 
4 1 2 18 20 
25 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
28 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 14 12 13 15 16 
14 1 2 3 4 9 9 9 9 9 9 9 9 18 9 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 12 14 15 13 16 
3 1 2 18 
24 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 16 14 12 13 15 16 
6 1 2 3 20 18 9 
4 1 2 18 20 
25 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 16 16 16 14 15 13 12 16 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
23 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
19 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 16 18 21 22 
26 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
54 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
4 1 2 18 20 
39 1 2 3 9 9 4 6 5 7 8 9 10 10 17 5 7 8 10 11 10 16 16 22 22 17 5 7 8 22 22 22 22 22 22 22 22 19 17 22 
3 1 2 18 
36 1 2 3 4 5 6 7 8 9 10 10 11 10 16 23 23 16 5 17 7 8 22 22 22 22 22 22 22 22 11 22 12 14 13 15 16 
12 1 2 3 20 9 9 9 9 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
29 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 16 22 14 13 15 12 16 
4 1 2 18 20 
3 1 2 18 
26 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 21 18 16 
26 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 22 16 16 16 22 16 14 15 12 13 16 
3 1 2 18 
3 1 2 18 
23 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
41 1 2 3 9 9 4 5 6 7 8 9 10 10 5 17 7 8 10 5 17 7 8 10 10 10 10 10 11 10 16 16 16 16 22 16 16 15 13 12 14 16 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 18 9 
35 1 2 20 3 20 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 16 22 22 22 16 16 14 15 13 12 16 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 20 18 20 
19 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 19 17 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 15 14 12 13 16 
37 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 5 17 7 8 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 17 19 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 18 21 16 
28 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 11 10 16 22 22 16 16 14 12 15 13 16 
3 1 2 18 
19 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
23 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 13 14 15 12 16 
3 1 2 18 
9 1 2 20 3 20 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
8 1 2 20 3 20 9 19 9 
22 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 18 21 22 
6 1 2 3 4 18 9 
4 1 2 18 20 
26 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
15 1 2 3 4 6 5 7 8 9 10 11 10 18 21 16 
36 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 16 16 16 16 16 16 22 22 14 12 13 15 16 
3 1 2 18 
17 1 2 3 20 4 6 5 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
34 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 11 10 16 16 14 15 13 12 16 
24 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 11 10 14 13 15 12 16 
32 1 2 3 4 6 5 7 8 9 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
20 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 15 14 12 13 16 
6 1 2 3 20 18 9 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
8 1 2 3 9 9 9 19 9 
28 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 16 22 14 12 13 15 16 
28 1 2 3 9 9 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 10 10 10 10 10 17 19 10 
24 1 2 20 3 20 4 6 5 7 8 9 5 17 7 8 10 10 11 10 14 13 12 15 16 
3 1 2 18 
6 1 2 20 20 18 20 
4 1 2 18 20 
3 1 2 18 
15 1 2 3 9 9 4 6 5 7 8 9 10 19 17 10 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
37 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
19 1 2 20 3 20 9 9 4 5 6 7 8 9 10 10 10 10 19 17 
25 1 2 3 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 19 17 10 
4 1 2 18 20 
19 1 2 3 4 6 5 7 8 9 10 10 10 11 10 12 13 15 14 16 
3 1 2 18 
24 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 13 15 12 14 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
26 1 2 3 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 11 10 12 13 15 14 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
27 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 14 13 12 15 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 20 4 5 6 7 8 9 10 11 10 14 13 15 12 16 
3 1 2 18 
24 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 23 16 22 15 13 12 14 22 
12 1 2 3 4 5 6 7 8 9 17 19 10 
43 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 17 5 7 8 10 10 10 10 10 17 19 10 
3 1 2 18 
57 1 2 3 20 9 9 4 6 5 7 8 9 5 17 7 8 10 5 17 7 8 10 10 10 17 5 7 8 10 10 10 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 22 16 22 22 14 12 15 13 16 
3 1 2 18 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 19 17 
3 1 2 18 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
30 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 11 10 16 16 22 22 22 22 22 22 12 14 13 15 16 
27 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
38 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
39 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 17 5 7 8 10 17 5 7 8 10 10 10 11 10 5 17 7 8 16 14 12 13 15 22 
31 1 2 20 3 20 9 4 6 5 7 8 9 10 5 17 7 8 10 17 5 7 8 10 10 10 10 10 10 10 19 17 
3 1 2 18 
31 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 16 16 16 22 22 22 16 13 14 15 12 16 
5 1 2 20 18 20 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
23 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 17 19 
18 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
24 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
28 1 2 20 3 20 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 16 14 12 13 15 16 
3 1 2 18 
26 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 14 13 12 15 16 
3 1 2 18 
6 1 2 3 4 18 9 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 21 18 16 
24 1 2 3 20 4 5 6 7 8 9 10 11 10 16 16 22 22 16 16 14 12 13 15 16 
4 1 2 18 20 
37 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 16 16 13 14 15 12 16 
15 1 2 3 4 6 5 7 8 9 10 11 10 21 18 16 
3 1 2 18 
5 1 2 3 18 9 
11 1 2 23 23 23 20 23 23 23 18 20 
19 1 2 3 4 5 6 7 8 9 11 10 16 16 16 14 12 15 13 16 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
16 1 2 3 4 6 5 7 8 9 11 10 14 12 15 13 16 
30 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
28 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 16 16 14 12 15 13 16 
3 1 2 18 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
18 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 17 19 10 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 15 13 14 12 16 
45 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 16 16 22 22 22 22 22 16 22 22 22 22 22 5 17 7 8 22 22 22 11 22 16 21 18 16 
29 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 17 19 10 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
14 1 2 3 4 6 5 7 8 9 10 10 18 21 10 
21 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 17 19 10 
3 1 2 18 
6 1 2 3 9 18 9 
3 1 2 18 
7 1 2 20 3 20 18 9 
4 1 2 18 20 
23 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 17 19 10 
19 1 2 3 20 4 5 6 7 8 9 10 11 10 16 14 12 13 15 16 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
9 1 2 3 9 9 9 9 9 19 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 17 19 10 
4 1 2 18 20 
18 1 2 3 20 4 5 6 7 8 9 10 11 10 15 14 13 12 16 
3 1 2 18 
7 1 2 3 9 9 19 9 
3 1 2 18 
27 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 14 12 15 13 16 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
6 1 2 3 20 18 9 
16 1 2 3 4 6 5 7 8 9 11 10 16 16 18 21 16 
64 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 22 22 22 22 16 22 22 22 5 17 7 8 16 15 12 14 13 22 
3 1 2 18 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 19 17 10 
5 1 2 20 18 20 
3 1 2 18 
6 1 2 20 20 18 20 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 14 13 12 15 16 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 13 15 12 16 
27 1 2 3 4 6 5 7 8 9 10 10 10 10 17 5 7 8 10 10 10 11 10 12 14 13 15 16 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 11 10 15 14 12 13 16 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 10 10 10 17 19 
17 1 2 3 20 4 6 5 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
5 1 2 3 19 9 
3 1 2 18 
19 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 19 17 10 
28 1 2 3 20 4 6 5 7 8 9 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
13 1 2 3 9 4 6 5 7 8 9 17 19 10 
22 1 2 3 4 9 5 6 7 8 9 5 17 7 8 10 10 10 10 10 19 17 10 
11 1 2 3 9 9 9 9 9 9 9 19 
3 1 2 18 
20 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 14 13 15 12 16 
28 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 22 16 16 16 16 16 22 22 15 14 13 12 22 
3 1 2 18 
39 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 11 10 16 16 22 22 22 22 16 16 17 5 7 8 16 15 13 12 14 22 
47 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 16 16 16 16 21 18 16 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
16 1 2 3 4 6 5 7 8 9 10 10 11 10 18 21 16 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 13 14 15 12 16 
4 1 2 18 20 
3 1 2 18 
37 1 2 3 20 9 4 6 5 7 8 9 5 17 7 8 10 17 5 7 8 10 17 5 7 8 10 5 17 7 8 10 10 10 10 19 17 10 
4 1 2 18 20 
27 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 17 19 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
9 1 2 20 3 20 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
8 1 2 3 20 9 4 19 9 
3 1 2 18 
24 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 17 5 7 8 10 10 19 17 10 
13 1 2 3 9 9 9 9 9 9 9 9 18 9 
26 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 14 13 12 15 16 
3 1 2 18 
20 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 19 17 10 
4 1 2 18 20 
22 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 17 19 10 
5 1 2 20 18 20 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
21 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 16 14 13 15 12 16 
38 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 22 16 16 13 12 14 15 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 10 10 11 10 21 18 16 
16 1 2 3 4 6 5 7 8 9 10 11 10 16 18 21 16 
6 1 2 3 9 19 9 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 11 10 14 15 13 12 16 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 3 19 9 
4 1 2 18 20 
29 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 5 17 7 8 10 10 10 10 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 9 18 9 
16 1 2 3 4 5 6 7 8 9 11 10 14 15 12 13 16 
6 1 2 3 20 18 9 
3 1 2 18 
10 1 2 20 20 3 20 9 9 18 9 
3 1 2 18 
24 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 14 13 15 12 16 
5 1 2 3 19 9 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
5 1 2 3 19 9 
5 1 2 20 18 20 
15 1 2 3 9 4 9 5 6 7 8 9 10 19 17 10 
3 1 2 18 
6 1 2 3 9 19 9 
4 1 2 18 20 
15 1 2 3 4 6 5 7 8 9 10 11 10 18 21 16 
16 1 2 3 9 9 9 4 5 6 7 8 9 10 19 17 10 
25 1 2 3 20 9 9 4 5 6 7 8 9 11 10 16 16 16 16 22 22 14 12 13 15 16 
28 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 22 22 22 22 22 14 13 12 15 16 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 19 17 10 
20 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 14 13 12 15 16 
32 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 11 10 21 18 16 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 14 12 13 15 16 
6 1 2 3 9 18 9 
3 1 2 18 
7 1 2 3 20 9 18 9 
15 1 2 3 20 4 6 5 7 8 9 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
24 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 16 14 12 13 15 16 
20 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 19 17 
4 1 2 18 20 
35 1 2 3 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 11 10 16 16 16 16 16 22 22 16 16 12 13 14 15 16 
29 1 2 3 9 4 5 6 7 8 9 10 11 10 16 5 17 7 8 22 22 22 22 11 22 13 12 14 15 16 
4 1 2 18 20 
9 1 2 3 20 9 9 9 18 9 
14 1 2 3 9 9 9 9 9 9 9 9 9 18 9 
28 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 23 16 16 22 21 18 22 
32 1 2 3 4 5 6 7 8 9 5 17 7 8 10 17 5 7 8 10 10 10 10 10 11 10 16 16 22 22 17 19 22 
27 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 14 13 15 12 16 
24 1 2 3 9 9 9 9 4 6 5 7 8 9 10 11 10 16 16 16 14 15 13 12 16 
11 1 2 3 20 9 9 9 9 9 19 9 
21 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 14 12 13 15 16 
39 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 16 16 16 22 22 22 22 22 22 22 16 5 17 7 8 16 13 15 12 14 22 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
24 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 22 22 22 22 22 22 17 19 22 
26 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 16 16 16 14 13 12 15 16 
7 1 2 3 20 9 19 9 
47 1 2 3 9 9 9 23 23 9 9 9 4 9 9 9 9 9 9 9 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 11 10 16 14 13 15 12 16 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 10 19 17 
29 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 13 14 15 12 16 
17 1 2 3 4 6 5 7 8 9 10 10 11 10 16 18 21 16 
25 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 11 10 16 16 16 18 21 16 
4 1 2 18 20 
30 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 11 10 18 21 16 
20 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 19 17 10 
5 1 2 3 18 9 
3 1 2 18 
23 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 16 16 14 12 15 13 16 
25 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 19 17 22 
3 1 2 18 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 21 18 16 
42 1 2 3 4 6 5 7 8 9 10 11 10 16 16 16 22 22 16 22 22 22 22 22 22 22 16 16 16 22 22 22 16 16 16 16 16 16 14 13 12 15 16 
19 1 2 3 4 5 6 7 8 9 11 10 16 22 22 14 13 12 15 16 
5 1 2 3 19 9 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
23 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 19 17 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 21 18 16 
24 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 19 17 10 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
63 1 2 3 20 4 6 5 7 8 9 11 10 16 22 16 16 22 22 22 22 22 17 5 7 8 22 22 22 22 22 22 22 22 11 22 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 13 14 12 15 16 
30 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 16 22 22 22 22 22 14 13 12 15 16 
6 1 2 3 20 18 9 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
3 1 2 18 
10 1 2 3 9 9 9 9 9 18 9 
33 1 2 20 3 20 9 9 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 19 17 
15 1 2 3 20 4 6 5 7 8 9 10 10 19 17 10 
5 1 2 20 18 20 
7 1 2 3 9 9 18 9 
25 1 2 3 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 10 10 11 10 21 18 16 
35 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 22 16 16 17 5 7 8 16 13 14 12 15 22 
26 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 16 14 13 12 15 16 
21 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 21 18 16 
7 1 2 20 3 20 18 9 
3 1 2 18 
5 1 2 20 18 20 
9 1 2 3 9 9 9 9 9 19 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
3 1 2 18 
8 1 2 3 9 9 9 18 9 
26 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 16 16 16 16 16 14 15 13 12 16 
23 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 16 16 14 13 15 12 16 
18 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 17 19 10 
20 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 11 10 21 18 16 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
19 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
88 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 11 22 16 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 17 19 22 
3 1 2 18 
4 1 2 18 20 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
33 1 2 3 4 6 5 7 8 9 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 12 14 15 13 16 
29 1 2 3 20 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 12 14 15 13 16 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
26 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
24 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
29 1 2 3 20 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 14 12 15 13 16 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
6 1 2 20 20 18 20 
3 1 2 18 
35 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
17 1 2 3 4 5 6 7 8 9 10 11 10 15 13 12 14 16 
22 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 13 14 15 12 16 
14 1 2 3 9 9 4 6 5 7 8 9 19 17 10 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
11 1 2 3 9 9 9 9 9 9 19 9 
3 1 2 18 
16 1 2 20 3 20 9 9 9 9 9 9 9 9 9 19 9 
23 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 15 14 12 13 16 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
22 1 2 3 20 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 17 19 10 
6 1 2 3 4 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
38 1 2 3 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 17 5 7 8 10 11 10 16 22 22 22 22 22 22 22 14 12 15 13 16 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 5 17 7 8 10 11 10 14 13 12 15 16 
21 1 2 3 4 6 5 7 8 9 5 17 7 8 10 11 10 12 13 15 14 16 
3 1 2 18 
15 1 2 3 20 4 6 5 7 8 9 10 10 21 18 10 
4 1 2 18 20 
21 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 16 13 14 12 15 16 
4 1 2 18 20 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 19 17 10 
23 1 2 3 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 17 19 10 
4 1 2 18 20 
18 1 2 3 20 9 9 4 6 5 7 8 9 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
30 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 16 16 16 16 22 22 22 16 16 16 14 15 13 12 16 
4 1 2 18 20 
13 1 2 3 9 4 6 5 7 8 9 17 19 10 
3 1 2 18 
32 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 5 17 7 8 10 10 10 10 10 11 10 13 12 15 14 16 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
15 1 2 3 4 6 5 7 8 9 10 10 10 17 19 10 
24 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 19 17 
23 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 18 21 10 
4 1 2 18 20 
13 1 2 3 9 4 6 5 7 8 9 19 17 10 
26 1 2 3 20 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 21 18 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
44 1 2 3 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 17 5 7 8 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 17 19 
21 1 2 3 20 4 5 6 7 8 9 10 17 5 7 8 10 10 10 19 17 10 
11 1 2 3 9 9 9 9 9 9 19 9 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
23 1 2 3 20 9 9 9 4 5 6 7 8 9 11 10 16 22 22 15 14 13 12 16 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
7 1 2 20 3 20 18 9 
36 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 5 17 7 8 10 5 17 7 8 10 10 10 11 10 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 20 18 9 
3 1 2 18 
5 1 2 3 19 9 
8 1 2 3 9 9 9 19 9 
5 1 2 3 18 9 
3 1 2 18 
7 1 2 3 20 9 18 9 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
22 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 11 10 14 13 12 15 16 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 14 12 13 15 16 
3 1 2 18 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
6 1 2 3 20 18 9 
23 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 17 19 
19 1 2 3 20 9 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
37 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 11 10 16 22 22 22 22 22 22 16 16 22 17 5 7 8 16 13 15 12 14 22 
4 1 2 18 20 
3 1 2 18 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
30 1 2 3 4 6 5 7 8 9 10 10 10 5 17 7 8 10 10 11 10 5 17 7 8 16 15 13 12 14 22 
26 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
17 1 2 3 4 5 6 7 8 9 10 11 10 16 16 18 21 22 
27 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 16 15 14 12 13 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
21 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
20 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 19 17 10 
4 1 2 18 20 
15 1 2 3 9 9 4 5 6 7 8 9 10 19 17 10 
16 1 2 3 20 9 9 4 5 6 7 8 9 10 10 17 19 
3 1 2 18 
10 1 2 3 9 9 9 9 9 9 19 
22 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 15 14 13 12 16 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 21 18 16 
14 1 2 3 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 4 19 9 
23 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
17 1 2 3 20 9 4 6 5 7 8 9 10 10 10 17 19 10 
3 1 2 18 
27 1 2 20 3 20 4 5 6 7 8 9 10 10 10 10 10 5 17 7 8 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
3 1 2 18 
24 1 2 3 9 4 6 5 7 8 9 11 10 16 16 23 16 16 16 16 15 13 12 14 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
46 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 16 16 16 22 22 22 22 22 22 16 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 13 14 15 12 22 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 12 14 13 15 16 
3 1 2 18 
21 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
5 1 2 3 19 9 
21 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 16 15 13 12 14 16 
24 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 14 12 15 13 16 
3 1 2 18 
42 1 2 3 20 9 4 6 5 7 8 9 10 10 17 5 7 8 10 10 10 11 10 16 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 21 18 16 
23 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 17 19 22 
3 1 2 18 
15 1 2 23 23 23 20 23 20 3 20 9 4 9 9 19 
3 1 2 18 
3 1 2 18 
24 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 14 15 12 13 22 
13 1 2 20 3 20 9 9 9 9 9 9 18 9 
12 1 2 3 4 5 6 7 8 9 18 21 10 
44 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 10 11 10 16 22 22 22 22 16 17 5 7 8 22 22 22 11 22 13 14 15 12 16 
16 1 2 3 20 4 5 6 7 8 9 10 10 10 21 18 10 
4 1 2 18 20 
33 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 11 10 16 22 22 22 22 12 13 15 14 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
51 1 2 3 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 5 17 7 8 10 10 17 5 7 8 10 5 17 7 8 10 10 17 5 7 8 10 10 10 11 10 16 16 14 15 12 13 16 
17 1 2 3 4 6 5 7 8 9 11 10 16 14 13 15 12 16 
31 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 11 10 16 16 22 22 22 22 22 14 13 15 12 16 
23 1 2 3 9 9 4 5 6 7 8 9 11 10 16 16 22 22 22 14 13 12 15 16 
16 1 2 3 9 9 4 5 6 7 8 9 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
5 1 2 3 18 9 
4 1 2 18 20 
20 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 11 10 18 21 16 
5 1 2 3 18 9 
25 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
3 1 2 18 
5 1 2 3 18 9 
36 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 16 16 22 17 5 7 8 22 22 22 22 14 15 13 12 22 
3 1 2 18 
23 1 2 3 9 9 9 9 4 6 5 7 8 9 11 10 16 22 22 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
31 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 17 5 7 8 22 22 22 22 11 22 16 13 14 15 12 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
14 1 2 3 4 6 5 7 8 9 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 10 19 17 
4 1 2 18 20 
20 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 13 14 15 12 16 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
3 1 2 18 
15 1 2 3 9 4 6 5 7 8 9 10 10 17 19 10 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
19 1 2 3 4 5 6 7 8 9 10 10 11 10 16 12 13 15 14 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 14 15 12 16 
7 1 2 3 9 4 18 9 
3 1 2 18 
21 1 2 3 9 9 9 9 4 9 6 5 7 8 9 10 10 11 10 18 21 16 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
9 1 2 3 9 9 9 9 19 9 
51 1 2 20 20 20 20 20 20 20 3 20 4 5 6 7 8 9 10 11 10 16 16 16 16 22 22 22 22 22 22 22 22 22 16 16 16 16 22 22 16 16 16 16 16 16 16 14 13 12 15 16 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 18 9 
18 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 19 17 
29 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 22 22 22 22 22 22 21 18 22 
5 1 2 3 19 9 
4 1 2 18 20 
8 1 2 3 9 9 9 18 9 
4 1 2 18 20 
6 1 2 3 20 18 9 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 14 13 15 12 16 
3 1 2 18 
26 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 22 22 22 22 22 22 22 17 19 22 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 12 13 15 16 
21 1 2 3 9 4 5 6 7 8 9 10 5 17 7 8 10 11 10 19 17 16 
16 1 2 3 4 6 5 7 8 9 11 10 12 13 15 14 16 
15 1 2 3 4 5 6 7 8 9 10 10 10 10 17 19 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
15 1 2 3 20 4 6 5 7 8 9 10 10 10 17 19 
19 1 2 3 9 9 4 5 6 7 8 9 10 11 10 14 13 15 12 16 
13 1 2 3 20 9 9 9 9 9 9 9 9 19 
30 1 2 20 3 20 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 17 5 7 8 16 13 14 12 15 22 
31 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 13 12 14 15 16 
3 1 2 18 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
20 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 16 21 18 16 
3 1 2 18 
35 1 2 20 20 20 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 5 17 7 8 10 10 11 10 16 22 14 12 13 15 16 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
27 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
31 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 16 16 16 16 22 22 16 22 22 22 17 19 22 
27 1 2 3 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 17 19 
32 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 17 19 10 
28 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 12 14 13 15 16 
4 1 2 18 20 
17 1 2 3 20 9 9 4 6 5 7 8 9 10 10 17 19 10 
16 1 2 3 20 4 6 5 7 8 9 10 10 10 19 17 10 
7 1 2 3 20 9 19 9 
7 1 2 3 20 9 9 19 
22 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 16 16 13 14 12 15 16 
28 1 2 20 3 20 4 6 5 7 8 9 10 10 10 11 10 16 16 16 23 16 16 16 13 14 12 15 16 
11 1 2 3 20 9 9 9 9 9 19 9 
6 1 2 3 20 18 9 
4 1 2 18 20 
22 1 2 20 20 3 20 4 6 5 7 8 9 10 11 10 16 16 14 12 13 15 16 
39 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
4 1 2 18 20 
6 1 2 20 20 18 20 
9 1 2 20 20 3 20 9 19 9 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
22 1 2 20 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
5 1 2 3 19 9 
3 1 2 18 
4 1 2 18 20 
30 1 2 3 20 4 5 6 7 8 9 10 11 10 16 16 23 16 16 16 16 22 22 22 22 22 12 14 15 13 16 
21 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 13 14 12 15 16 
4 1 2 18 20 
29 1 2 20 3 20 9 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 10 11 10 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 15 13 12 14 16 
4 1 2 18 20 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
12 1 2 3 4 5 6 7 8 9 17 19 10 
3 1 2 18 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
7 1 2 3 20 9 18 9 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 9 18 9 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 15 14 13 12 16 
4 1 2 18 20 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
3 1 2 18 
23 1 2 20 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 19 
7 1 2 3 20 9 18 9 
21 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 18 21 16 
18 1 2 3 9 4 5 6 7 8 9 11 10 16 13 14 12 15 16 
23 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 11 10 16 14 13 12 15 16 
3 1 2 18 
26 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 11 10 16 16 16 13 14 12 15 16 
25 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 16 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
18 1 2 3 9 9 4 5 6 7 8 9 11 10 13 15 12 14 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
23 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 14 15 13 12 16 
10 1 2 3 20 9 9 9 9 18 9 
4 1 2 18 20 
32 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 11 10 16 23 23 23 23 16 22 22 22 22 14 13 15 12 16 
3 1 2 18 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
22 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 13 14 12 15 16 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 18 9 
19 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 17 19 10 
16 1 2 3 20 4 6 5 7 8 9 10 10 10 10 19 17 
12 1 2 3 4 5 6 7 8 9 19 17 10 
12 1 2 3 20 9 9 9 9 9 9 18 9 
40 1 2 3 4 6 5 7 8 9 10 11 10 16 16 16 16 22 22 16 16 22 22 17 5 7 8 22 22 22 22 22 22 11 22 16 14 13 12 15 16 
5 1 2 3 18 9 
5 1 2 20 18 20 
32 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 14 13 12 15 16 
3 1 2 18 
6 1 2 3 20 18 9 
12 1 2 3 20 9 9 9 9 9 9 18 9 
22 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 22 14 12 13 15 16 
29 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
32 1 2 3 20 9 9 4 6 5 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 16 16 12 14 13 15 16 
19 1 2 3 9 9 4 6 5 7 8 9 11 10 16 14 12 15 13 16 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
16 1 2 3 20 4 5 6 7 8 9 11 10 16 21 18 16 
4 1 2 18 20 
37 1 2 3 20 4 6 5 7 8 9 11 10 16 23 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 13 14 15 12 16 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
11 1 2 20 3 20 9 9 9 9 19 9 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
48 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 5 17 7 8 22 14 13 15 12 22 
19 1 2 20 3 20 4 5 6 7 8 9 10 11 10 14 13 12 15 16 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
31 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 11 10 13 12 14 15 16 
3 1 2 18 
33 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 16 22 22 22 16 16 22 22 16 16 22 22 14 13 15 12 16 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
5 1 2 20 18 20 
16 1 2 3 4 6 5 7 8 9 11 10 13 14 12 15 16 
3 1 2 18 
8 1 2 3 20 9 9 19 9 
3 1 2 18 
26 1 2 3 4 5 6 7 8 9 11 10 16 22 22 16 16 16 22 22 16 16 13 12 15 14 16 
5 1 2 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
17 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 19 17 
40 1 2 20 3 20 9 4 6 5 7 8 9 10 17 5 7 8 10 5 17 7 8 10 10 5 17 7 8 10 10 11 10 16 22 22 13 14 15 12 16 
23 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 22 22 13 14 15 12 16 
53 1 2 3 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 10 10 11 10 16 16 16 16 17 5 7 8 22 22 22 22 11 22 16 16 12 13 15 14 16 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 12 13 15 14 16 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 13 12 14 15 16 
3 1 2 18 
3 1 2 18 
39 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 16 16 16 16 16 22 5 17 7 8 22 22 22 11 22 16 16 16 22 14 13 12 15 16 
29 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 16 22 22 16 22 22 22 16 12 14 13 15 16 
4 1 2 18 20 
6 1 2 3 20 19 9 
36 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 16 16 16 22 22 22 16 22 22 22 22 16 16 13 14 12 15 16 
8 1 2 3 20 9 9 19 9 
22 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 11 10 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
19 1 2 3 9 9 4 5 6 7 8 9 11 10 16 14 12 13 15 16 
15 1 2 3 20 4 6 5 7 8 9 10 10 10 17 19 
16 1 2 3 9 9 9 4 6 5 7 8 9 10 19 17 10 
31 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 18 21 16 
4 1 2 18 20 
30 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 17 19 
36 1 2 3 4 6 5 7 8 9 10 11 10 16 16 22 22 22 22 22 16 22 22 5 17 7 8 22 22 22 11 22 13 14 12 15 16 
4 1 2 18 20 
10 1 2 3 9 9 9 9 9 9 19 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 14 13 12 15 16 
5 1 2 20 18 20 
4 1 2 18 20 
43 1 2 3 20 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 11 10 16 22 22 16 14 12 13 15 16 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 19 
32 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 14 13 15 12 16 
7 1 2 3 20 9 18 9 
3 1 2 18 
8 1 2 3 9 9 9 19 9 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 18 9 
6 1 2 3 20 19 9 
3 1 2 18 
40 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 16 16 16 16 16 5 17 7 8 22 22 22 22 11 22 16 22 22 22 14 12 13 15 16 
5 1 2 3 18 9 
20 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 19 17 
53 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 5 17 7 8 10 17 5 7 8 10 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 16 22 22 22 14 15 12 13 22 
32 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 16 16 22 22 22 16 22 22 22 22 22 22 18 21 22 
3 1 2 18 
33 1 2 3 4 6 5 7 8 9 10 10 17 5 7 8 10 10 11 10 16 16 22 22 22 22 22 22 22 14 12 13 15 16 
60 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 5 17 7 8 10 17 5 7 8 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 17 5 7 8 16 11 22 14 12 15 13 16 
3 1 2 18 
7 1 2 3 9 9 18 9 
35 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 17 5 7 8 10 17 5 7 8 10 10 10 10 11 10 13 14 12 15 16 
4 1 2 18 20 
9 1 2 3 20 9 9 9 19 9 
48 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 11 22 15 13 12 14 16 
3 1 2 18 
3 1 2 18 
20 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 13 14 12 15 16 
6 1 2 3 20 18 9 
27 1 2 3 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 10 17 19 
40 1 2 3 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 5 17 7 8 10 17 5 7 8 10 10 10 11 10 16 22 22 15 13 12 14 16 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 19 17 10 
23 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 12 13 15 14 16 
3 1 2 18 
14 1 2 3 9 4 5 6 7 8 9 10 19 17 10 
5 1 2 20 18 20 
23 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
36 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 5 17 7 8 10 10 11 10 16 22 22 22 22 16 22 22 14 15 13 12 22 
5 1 2 3 18 9 
9 1 2 20 3 20 9 9 18 9 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
5 1 2 3 19 9 
5 1 2 20 18 20 
38 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 21 18 16 
3 1 2 18 
15 1 2 3 4 6 5 7 8 9 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
10 1 2 3 20 9 9 9 9 9 19 
17 1 2 3 9 4 6 5 7 8 9 10 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
6 1 2 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
29 1 2 3 4 6 5 7 8 9 5 17 7 8 10 11 10 16 16 16 5 17 7 8 16 13 14 15 12 22 
23 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
3 1 2 18 
15 1 2 3 20 9 4 6 5 7 8 9 10 19 17 10 
22 1 2 20 3 20 9 4 6 5 7 8 9 11 10 16 22 22 14 12 15 13 16 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
8 1 2 3 9 9 9 19 9 
3 1 2 18 
46 1 2 3 9 9 4 5 6 7 8 9 11 10 16 23 16 22 22 17 5 7 8 22 22 22 22 11 22 16 22 22 22 22 22 22 22 22 22 22 22 16 13 15 12 14 16 
24 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 19 17 
35 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 5 17 7 8 10 5 17 7 8 10 10 10 10 17 19 10 
3 1 2 18 
15 1 2 3 20 4 6 5 7 8 9 10 10 18 21 10 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
16 1 2 3 20 9 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
7 1 2 3 9 9 18 9 
17 1 2 3 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
5 1 2 23 18 23 
26 1 2 3 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 5 17 7 8 10 19 17 10 
5 1 2 3 18 9 
4 1 2 18 20 
9 1 2 3 9 9 9 9 9 19 
3 1 2 18 
8 1 2 20 20 20 20 18 20 
5 1 2 20 18 20 
5 1 2 20 18 20 
49 1 2 20 3 20 9 9 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 10 17 5 7 8 10 10 5 17 7 8 10 17 5 7 8 10 10 10 11 10 14 15 12 13 16 
21 1 2 3 20 9 4 6 5 7 8 9 5 17 7 8 10 11 10 21 18 16 
34 1 2 3 20 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 16 22 22 22 16 17 5 7 8 22 22 22 17 19 22 
6 1 2 3 20 19 9 
6 1 2 3 20 19 9 
23 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 19 17 
39 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 5 17 7 8 10 10 11 10 16 17 5 7 8 16 14 12 13 15 22 
38 1 2 3 20 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
28 1 2 20 20 20 20 20 20 20 3 20 9 9 4 5 6 7 8 9 11 10 16 16 12 14 13 15 16 
4 1 2 18 20 
6 1 2 3 20 18 9 
9 1 2 3 20 9 9 9 19 9 
30 1 2 3 20 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
41 1 2 3 20 4 6 5 7 8 9 11 10 16 16 16 16 16 16 16 16 16 16 16 16 16 22 22 22 22 22 22 22 22 22 22 22 14 15 12 13 16 
33 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 16 16 22 22 22 5 17 7 8 22 22 22 17 19 22 
3 1 2 18 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 10 11 10 16 13 12 14 15 16 
46 1 2 3 9 4 6 5 7 8 9 11 10 17 5 7 8 16 22 22 22 22 22 22 22 22 22 22 17 5 7 8 22 22 11 22 16 16 16 16 16 16 13 14 12 15 16 
4 1 2 18 20 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
29 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
24 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 17 19 10 
27 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
7 1 2 3 9 9 9 19 
19 1 2 3 9 9 9 4 5 6 7 8 9 11 10 14 12 15 13 16 
4 1 2 18 20 
31 1 2 3 9 4 6 5 7 8 9 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 11 10 16 21 18 16 
18 1 2 3 4 6 5 7 8 9 11 10 16 23 12 13 14 15 16 
3 1 2 18 
7 1 2 3 9 9 18 9 
46 1 2 3 20 9 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 22 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 17 19 22 
12 1 2 3 4 6 5 7 8 9 19 17 10 
3 1 2 18 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
17 1 2 3 9 9 4 5 6 7 8 9 11 10 16 18 21 16 
17 1 2 3 9 4 6 5 7 8 9 11 10 14 12 13 15 16 
27 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 19 17 
24 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 11 10 16 22 18 21 22 
3 1 2 18 
7 1 2 3 9 9 19 9 
3 1 2 18 
3 1 2 18 
20 1 2 3 20 9 4 6 5 7 8 9 10 10 11 10 13 14 12 15 16 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 13 15 12 16 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
27 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 11 10 16 16 22 12 13 15 14 16 
30 1 2 3 20 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 10 10 10 10 11 10 16 16 21 18 16 
22 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 13 14 15 12 16 
21 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 17 19 10 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 18 21 16 
44 1 2 3 20 4 6 5 7 8 9 5 17 7 8 10 10 17 5 7 8 10 17 5 7 8 10 10 17 5 7 8 10 10 10 10 10 11 10 16 12 15 13 14 16 
4 1 2 18 20 
13 1 2 3 20 9 9 9 9 9 9 9 19 9 
24 1 2 3 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
5 1 2 23 18 23 
33 1 2 3 20 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 21 18 22 
3 1 2 18 
3 1 2 18 
31 1 2 3 20 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 17 19 
15 1 2 3 4 6 5 7 8 9 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
8 1 2 20 3 20 9 18 9 
3 1 2 18 
25 1 2 3 9 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 14 12 13 15 16 
33 1 2 3 4 5 6 7 8 9 5 17 7 8 10 11 10 16 22 22 22 22 22 16 16 16 22 22 22 16 16 21 18 16 
4 1 2 18 20 
12 1 2 20 3 20 9 9 9 9 9 9 19 
37 1 2 3 20 9 4 5 6 7 8 9 10 11 10 5 17 7 8 16 22 22 22 22 17 5 7 8 22 22 22 11 22 15 14 12 13 16 
3 1 2 18 
17 1 2 3 9 4 5 6 7 8 9 11 10 13 12 14 15 16 
30 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 22 22 18 21 22 
3 1 2 18 
18 1 2 3 9 9 9 9 4 5 6 7 8 9 11 10 18 21 16 
34 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 18 21 10 
5 1 2 3 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 17 19 16 
10 1 2 20 20 20 20 20 20 18 20 
4 1 2 18 20 
27 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
14 1 2 3 4 5 6 7 8 9 11 10 21 18 16 
3 1 2 18 
4 1 2 18 20 
30 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 22 22 15 13 12 14 16 
7 1 2 3 20 9 18 9 
8 1 2 3 9 9 9 18 9 
3 1 2 18 
33 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 16 16 22 22 22 22 22 22 16 14 13 15 12 16 
4 1 2 18 20 
41 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
46 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
30 1 2 3 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 10 10 11 10 16 16 22 14 13 12 15 16 
13 1 2 23 23 20 23 3 20 9 9 9 9 19 
3 1 2 18 
14 1 2 3 20 4 5 6 7 8 9 10 21 18 10 
3 1 2 18 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
22 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
8 1 2 3 20 9 9 9 19 
3 1 2 18 
9 1 2 23 23 23 20 23 18 20 
44 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
22 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 19 17 10 
15 1 2 3 4 6 5 7 8 9 10 10 10 17 19 10 
8 1 2 3 9 9 9 19 9 
27 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
31 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 19 17 
17 1 2 3 9 4 5 6 7 8 9 11 10 13 15 12 14 16 
14 1 2 3 4 6 5 7 8 9 11 10 18 21 16 
21 1 2 20 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 19 17 10 
21 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 11 10 21 18 16 
6 1 2 3 20 18 9 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 18 21 16 
4 1 2 18 20 
3 1 2 18 
45 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 16 16 16 16 22 22 17 5 7 8 22 22 22 22 22 22 22 11 22 16 14 15 13 12 16 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 19 9 
35 1 2 3 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 11 10 16 16 16 22 22 22 22 22 16 16 12 14 13 15 16 
3 1 2 18 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 17 19 10 
5 1 2 3 19 9 
31 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 14 12 13 15 16 
18 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 19 17 10 
20 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 18 21 16 
3 1 2 18 
23 1 2 3 9 9 4 5 6 7 8 9 11 10 16 16 16 22 22 12 15 13 14 16 
7 1 2 3 9 9 18 9 
7 1 2 3 9 9 19 9 
3 1 2 18 
33 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
21 1 2 3 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 21 18 10 
5 1 2 3 18 9 
3 1 2 18 
16 1 2 3 20 4 6 5 7 8 9 10 11 10 18 21 16 
21 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
11 1 2 3 20 9 9 9 9 9 19 9 
7 1 2 20 20 20 18 20 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 10 19 17 
8 1 2 3 9 9 9 19 9 
39 1 2 3 9 9 9 9 4 6 5 7 8 9 11 10 16 16 22 22 5 17 7 8 22 22 22 5 17 7 8 22 22 11 22 14 15 13 12 16 
3 1 2 18 
19 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 17 19 10 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
20 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 10 19 
19 1 2 3 4 6 5 7 8 9 10 11 10 16 16 22 22 18 21 22 
4 1 2 18 20 
5 1 2 3 19 9 
4 1 2 18 20 
4 1 2 18 20 
27 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 21 18 16 
4 1 2 18 20 
39 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 12 15 14 13 16 
3 1 2 18 
4 1 2 18 20 
23 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 14 13 12 15 16 
27 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
16 1 2 3 4 5 6 7 8 9 11 10 14 13 12 15 16 
29 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 16 22 22 22 22 16 17 19 22 
31 1 2 3 20 4 5 6 7 8 9 10 17 5 7 8 10 17 5 7 8 10 10 10 11 10 16 16 16 21 18 16 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
36 1 2 3 9 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 
8 1 2 3 9 9 9 9 19 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 21 18 16 
21 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 22 12 15 14 13 16 
3 1 2 18 
20 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 16 16 21 18 16 
27 1 2 20 3 20 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 16 16 14 12 13 15 16 
21 1 2 3 4 5 6 7 8 9 11 10 16 16 16 16 16 13 15 12 14 16 
5 1 2 20 18 20 
22 1 2 3 20 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 17 19 10 
29 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 22 22 16 13 14 15 12 16 
9 1 2 3 20 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 23 18 23 
25 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 14 13 12 15 16 
9 1 2 20 20 3 20 9 18 9 
18 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 17 19 10 
18 1 2 20 20 20 20 20 3 20 4 5 6 7 8 9 19 17 10 
30 1 2 20 20 3 20 9 4 6 5 7 8 9 10 9 9 9 9 9 9 9 9 9 9 9 9 10 19 17 10 
5 1 2 20 18 20 
3 1 2 18 
20 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 14 12 13 15 16 
20 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 19 17 
25 1 2 3 20 4 6 5 7 8 9 10 17 5 7 8 10 11 10 16 16 14 15 13 12 16 
37 1 2 20 20 20 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 16 5 17 7 8 16 14 12 13 15 22 
5 1 2 3 19 9 
3 1 2 18 
4 1 2 18 20 
23 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
46 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 18 21 16 
30 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 17 5 7 8 10 11 10 16 16 16 15 13 12 14 16 
3 1 2 18 
4 1 2 18 20 
8 1 2 20 3 20 4 19 9 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 18 21 16 
5 1 2 3 18 9 
3 1 2 18 
6 1 2 20 20 18 20 
22 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
6 1 2 3 9 19 9 
3 1 2 18 
6 1 2 3 9 18 9 
9 1 2 3 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
25 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
34 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 5 17 7 8 10 10 10 11 10 17 5 7 8 16 14 13 12 15 22 
15 1 2 20 20 3 20 9 9 9 9 9 9 9 19 9 
30 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 16 16 16 16 16 16 22 22 22 16 14 13 12 15 16 
4 1 2 18 20 
8 1 2 3 9 9 9 18 9 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 10 10 11 10 16 18 21 16 
33 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 17 19 
22 1 2 3 20 9 9 4 6 5 7 8 9 11 10 16 22 22 15 14 12 13 16 
4 1 2 18 20 
25 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 11 10 13 14 15 12 16 
8 1 2 20 3 20 9 18 9 
9 1 2 20 20 20 3 20 19 9 
39 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 16 14 12 15 13 16 
13 1 2 3 20 9 9 9 9 9 9 9 19 9 
3 1 2 18 
25 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
10 1 2 3 9 9 9 9 9 9 19 
47 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 17 5 7 8 10 10 17 5 7 8 10 10 10 11 10 16 16 16 16 22 22 16 5 17 7 8 16 14 12 13 15 22 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
36 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 16 16 22 22 22 22 22 22 17 5 7 8 22 22 17 19 22 
3 1 2 18 
5 1 2 3 18 9 
17 1 2 3 9 4 6 5 7 8 9 11 10 14 13 15 12 16 
6 1 2 3 20 18 9 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 19 
4 1 2 18 20 
27 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 13 14 15 12 16 
10 1 2 20 3 20 9 9 9 18 9 
3 1 2 18 
6 1 2 3 20 18 9 
14 1 2 3 20 9 9 9 9 9 9 9 9 18 9 
26 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 5 17 7 8 10 10 19 17 10 
27 1 2 20 3 20 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 16 12 13 15 14 16 
41 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 16 16 16 16 16 16 22 16 22 22 22 17 5 7 8 22 22 11 22 13 14 12 15 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
63 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 5 17 7 8 10 10 10 11 10 16 16 22 22 22 22 22 16 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 16 16 22 22 22 22 22 16 14 15 12 13 16 
4 1 2 18 20 
38 1 2 20 20 20 20 3 20 9 9 4 6 5 7 8 9 17 5 7 8 10 10 17 5 7 8 10 10 10 10 11 10 16 14 12 15 13 16 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 12 15 13 14 16 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
11 1 2 3 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
10 1 2 20 20 20 20 20 20 18 20 
6 1 2 3 9 19 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
25 1 2 3 20 9 9 4 5 6 7 8 9 11 10 16 22 22 22 16 16 15 12 13 14 16 
3 1 2 18 
16 1 2 3 20 4 6 5 7 8 9 10 11 10 21 18 16 
10 1 2 3 20 9 9 9 9 19 9 
6 1 2 20 23 18 23 
6 1 2 3 20 18 9 
5 1 2 20 18 20 
14 1 2 3 20 4 5 6 7 8 9 10 17 19 10 
42 1 2 20 20 3 20 9 9 9 9 4 5 6 7 8 9 11 10 16 16 16 16 22 22 22 17 5 7 8 22 22 22 22 22 11 22 16 12 13 15 14 16 
27 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
9 1 2 20 3 20 9 9 18 9 
28 1 2 3 4 5 6 7 8 9 11 10 16 16 16 22 22 22 22 16 16 22 22 16 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 18 9 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 14 13 15 12 16 
8 1 2 3 9 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
8 1 2 20 3 20 9 18 9 
7 1 2 3 20 9 18 9 
27 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 22 14 12 13 15 16 
15 1 2 3 4 5 6 7 8 9 10 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
41 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 5 17 7 8 10 5 17 7 8 10 10 11 10 16 16 16 5 17 7 8 16 14 13 15 12 22 
7 1 2 3 9 9 19 9 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 18 21 16 
52 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 10 17 5 7 8 10 10 10 10 11 10 16 16 16 16 22 22 22 22 22 22 22 17 5 7 8 16 13 14 12 15 22 
3 1 2 18 
6 1 2 3 9 18 9 
10 1 2 3 9 9 9 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 20 18 20 
5 1 2 20 18 20 
22 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
11 1 2 3 9 9 9 9 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
42 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 17 5 7 8 10 17 5 7 8 10 11 10 16 22 22 22 22 16 13 14 12 15 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
31 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 16 16 16 16 16 16 22 22 16 16 13 12 15 14 16 
11 1 2 20 3 20 9 9 9 9 18 9 
3 1 2 18 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
4 1 2 18 20 
26 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 20 18 20 
18 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 17 19 10 
14 1 2 3 4 6 5 7 8 9 11 10 21 18 16 
3 1 2 18 
4 1 2 18 20 
27 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
22 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 18 21 16 
4 1 2 18 20 
5 1 2 20 18 20 
25 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 13 15 12 14 16 
3 1 2 18 
7 1 2 3 20 4 18 9 
3 1 2 18 
17 1 2 3 9 4 6 5 7 8 9 10 10 11 10 18 21 16 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 9 19 9 
32 1 2 3 4 6 5 7 8 9 10 10 5 17 7 8 10 10 10 5 17 7 8 10 10 10 10 5 17 7 8 10 10 
7 1 2 3 20 9 18 9 
3 1 2 18 
41 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 11 10 16 14 15 13 12 16 
12 1 2 3 4 5 6 7 8 9 17 19 10 
4 1 2 18 20 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 9 9 9 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
10 1 2 3 9 9 9 9 9 9 19 
16 1 2 3 9 9 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
13 1 2 3 4 5 6 7 8 9 10 18 21 10 
7 1 2 3 9 9 18 9 
19 1 2 3 20 4 5 6 7 8 9 10 11 10 16 12 14 15 13 16 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
20 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 13 14 12 15 16 
4 1 2 18 20 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
5 1 2 20 18 20 
3 1 2 18 
23 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 14 13 12 15 16 
4 1 2 18 20 
22 1 2 3 4 5 6 7 8 9 17 5 7 8 10 11 10 16 13 14 15 12 16 
5 1 2 20 18 20 
53 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 17 5 7 8 10 5 17 7 8 10 10 10 5 17 7 8 10 17 5 7 8 10 10 10 11 10 5 17 7 8 16 13 15 14 12 22 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
39 1 2 3 20 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 11 10 16 16 22 22 5 17 7 8 16 14 15 13 12 22 
23 1 2 3 9 9 9 9 4 6 5 7 8 9 11 10 16 16 22 13 14 15 12 16 
18 1 2 3 20 9 4 6 5 7 8 9 10 11 10 16 21 18 22 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
26 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 21 18 10 
3 1 2 18 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
43 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 16 16 22 22 22 22 22 15 14 12 13 16 
46 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 17 5 7 8 10 17 5 7 8 10 10 17 5 7 8 10 10 11 10 16 22 22 22 22 22 22 13 14 15 12 16 
4 1 2 18 20 
30 1 2 3 20 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 16 22 22 22 22 12 13 15 14 16 
21 1 2 3 20 4 6 5 7 8 9 10 11 10 16 16 16 14 12 15 13 16 
3 1 2 18 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
39 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 5 17 7 8 10 10 10 10 11 10 18 21 16 
46 1 2 3 20 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 5 17 7 8 16 22 22 22 22 22 22 22 22 22 22 22 22 11 22 15 13 12 14 16 
20 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 13 14 15 12 16 
3 1 2 18 
4 1 2 18 20 
31 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 5 17 7 8 22 22 22 11 22 13 14 12 15 16 
3 1 2 18 
18 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
27 1 2 3 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
82 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 16 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 12 14 13 15 22 
45 1 2 3 9 4 5 6 7 8 9 11 10 16 16 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
42 1 2 3 9 4 6 5 7 8 9 11 10 16 16 22 22 22 22 22 22 5 17 7 8 22 17 5 7 8 22 22 22 22 22 22 11 22 14 13 12 15 16 
82 1 2 3 4 5 6 7 8 9 5 17 7 8 10 11 10 16 5 17 7 8 16 22 22 22 17 5 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 16 22 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 22 22 22 22 22 22 17 19 22 
3 1 2 18 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
57 1 2 3 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 17 5 7 8 10 10 11 10 16 16 22 22 22 16 22 22 22 22 22 22 16 16 22 22 22 22 22 22 22 22 14 15 13 12 16 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 12 15 13 14 16 
38 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 19 17 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
21 1 2 3 4 6 5 7 8 9 10 10 10 17 5 7 8 10 10 19 17 10 
5 1 2 20 18 20 
20 1 2 3 9 9 9 9 4 6 5 7 8 9 11 10 13 14 15 12 16 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
34 1 2 3 20 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
24 1 2 3 4 5 6 7 8 9 11 10 16 16 16 12 15 13 16 16 16 16 16 16 16 
33 1 2 3 9 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 22 16 14 12 13 15 16 
6 1 2 3 20 18 9 
4 1 2 18 20 
40 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 19 17 16 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
27 1 2 3 4 5 6 7 8 9 11 10 16 16 16 16 16 22 22 22 16 16 16 15 12 14 13 16 
3 1 2 18 
3 1 2 18 
18 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 19 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
4 1 2 18 20 
21 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 22 14 13 12 15 22 
13 1 2 3 20 4 6 5 7 8 9 17 19 10 
32 1 2 3 20 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 11 10 16 16 22 22 22 22 12 14 13 15 16 
3 1 2 18 
3 1 2 18 
8 1 2 20 3 20 9 18 9 
5 1 2 20 18 20 
20 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
29 1 2 20 20 20 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
6 1 2 20 20 18 20 
7 1 2 20 3 20 19 9 
7 1 2 3 9 4 19 9 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
21 1 2 3 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 18 21 10 
19 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 17 19 10 
3 1 2 18 
5 1 2 20 18 20 
25 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
5 1 2 20 18 20 
22 1 2 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 17 19 16 
32 1 2 3 20 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
16 1 2 20 3 20 4 6 5 7 8 9 10 10 10 17 19 
5 1 2 20 18 20 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
8 1 2 3 20 9 9 18 9 
5 1 2 20 18 20 
5 1 2 20 18 20 
7 1 2 20 3 20 18 9 
4 1 2 18 20 
15 1 2 3 20 9 4 6 5 7 8 9 10 19 17 10 
22 1 2 3 20 4 5 6 7 8 9 11 10 16 16 16 22 22 15 13 12 14 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
4 1 2 18 20 
26 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 14 13 12 15 16 
13 1 2 3 20 9 9 9 9 9 9 9 19 9 
24 1 2 3 20 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 14 12 15 13 16 
24 1 2 3 20 9 4 5 6 7 8 9 11 10 16 16 22 22 22 22 13 14 15 12 16 
22 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 19 17 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
36 1 2 3 20 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 11 10 16 16 16 16 16 16 16 22 16 16 13 14 12 15 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
26 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 16 22 22 22 22 22 22 19 17 22 
3 1 2 18 
9 1 2 3 20 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 18 9 
24 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 16 16 14 12 15 13 16 
6 1 2 3 20 18 9 
5 1 2 3 18 9 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 20 9 18 9 
48 1 2 3 4 6 5 7 8 9 11 10 16 5 17 7 8 16 11 22 17 5 7 8 16 22 22 22 22 17 5 7 8 22 22 22 22 22 11 22 16 22 22 22 14 15 12 13 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
8 1 2 3 9 9 9 19 9 
20 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 17 19 10 
7 1 2 3 20 9 18 9 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 11 10 13 12 14 15 16 
19 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 21 18 16 
29 1 2 3 9 4 5 6 7 8 9 10 5 17 7 8 10 10 11 10 5 17 7 8 16 13 14 12 15 22 
4 1 2 18 20 
3 1 2 18 
23 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 12 13 15 14 16 
47 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 17 5 7 8 10 10 11 10 16 16 22 22 22 22 22 22 22 22 16 22 22 22 16 16 22 22 22 22 18 21 16 
29 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
4 1 2 18 20 
28 1 2 3 20 9 4 6 5 7 8 9 10 10 10 17 5 7 8 10 10 11 10 16 16 16 18 21 16 
3 1 2 18 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 19 17 10 
28 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 16 16 22 22 22 22 22 14 15 13 12 16 
3 1 2 18 
6 1 2 3 20 18 9 
44 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 11 10 16 16 16 16 22 22 22 22 22 22 13 15 12 14 16 
31 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 14 13 15 12 16 
20 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 14 12 13 15 16 
49 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 16 16 16 16 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 13 15 12 14 16 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
40 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 22 16 16 22 22 22 22 22 22 22 22 22 22 22 16 16 14 15 12 13 16 
6 1 2 3 9 18 9 
15 1 2 3 9 4 6 5 7 8 9 11 10 18 21 16 
50 1 2 3 20 9 4 5 6 7 8 9 10 17 5 7 8 10 5 17 7 8 10 10 10 10 10 10 11 10 16 16 16 16 16 22 16 22 22 16 16 17 5 7 8 16 14 15 13 12 22 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
23 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 14 13 15 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 17 19 10 
27 1 2 3 20 4 5 6 7 8 9 10 11 10 16 16 16 16 22 22 22 22 16 13 14 12 15 16 
19 1 2 3 4 6 5 7 8 9 11 10 16 16 16 14 12 13 15 16 
29 1 2 3 20 9 4 5 6 7 8 9 11 10 16 16 17 5 7 8 16 22 22 11 22 15 13 12 14 16 
16 1 2 3 20 4 6 5 7 8 9 10 10 10 17 19 10 
27 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 17 5 7 8 10 10 11 10 16 18 21 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 4 19 9 
3 1 2 18 
29 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 5 17 7 8 16 14 12 15 13 22 
7 1 2 3 9 9 19 9 
27 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 16 22 22 22 22 22 16 15 12 14 13 16 
3 1 2 18 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
15 1 2 3 9 9 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
3 1 2 18 
19 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 19 17 10 
21 1 2 3 4 6 5 7 8 9 11 10 16 22 22 16 16 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 22 22 12 14 13 15 16 
4 1 2 18 20 
4 1 2 18 20 
24 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
6 1 2 20 20 18 20 
26 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 16 16 14 12 13 15 16 
5 1 2 3 19 9 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 14 15 12 16 
5 1 2 23 18 23 
3 1 2 18 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 15 13 12 14 16 
10 1 2 3 9 9 9 9 4 19 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
15 1 2 3 4 6 5 7 8 9 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
17 1 2 3 20 4 5 6 7 8 9 11 10 12 13 15 14 16 
3 1 2 18 
30 1 2 3 9 4 6 5 7 8 9 10 10 5 17 7 8 10 10 11 10 16 22 22 16 22 22 22 19 17 22 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
10 1 2 20 3 20 9 9 9 9 19 
25 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 9 18 9 
24 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 14 13 12 15 16 
9 1 2 20 3 20 9 9 19 9 
3 1 2 18 
44 1 2 3 20 9 9 4 6 5 7 8 9 10 10 17 5 7 8 10 5 17 7 8 10 17 5 7 8 10 5 17 7 8 10 10 11 10 16 22 22 22 17 19 22 
7 1 2 3 20 9 18 9 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
25 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
29 1 2 3 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 11 10 14 12 13 15 16 
18 1 2 3 9 4 6 5 7 8 9 11 10 16 13 12 14 15 16 
10 1 2 3 20 9 9 9 9 18 9 
8 1 2 3 9 9 9 18 9 
29 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 16 14 13 15 12 16 
27 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 16 22 22 22 22 22 22 16 16 18 21 16 
4 1 2 18 20 
11 1 2 3 20 9 9 9 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
8 1 2 3 9 9 9 19 9 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
27 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 11 10 14 12 13 15 16 
11 1 2 3 9 9 9 9 9 9 19 9 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
22 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
23 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
30 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 16 16 16 16 16 14 13 15 12 16 
15 1 2 3 4 5 6 7 8 9 10 11 10 18 21 16 
4 1 2 18 20 
3 1 2 18 
24 1 2 3 20 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 14 13 12 15 16 
10 1 2 3 20 9 9 9 9 9 19 
3 1 2 18 
11 1 2 20 20 3 20 9 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
29 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 17 5 7 8 10 10 
7 1 2 3 9 9 18 9 
30 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 5 17 7 8 10 11 10 16 14 13 12 15 16 
4 1 2 18 20 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
50 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 16 16 16 13 14 15 12 16 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 18 21 16 
3 1 2 18 
5 1 2 3 18 9 
3 1 2 18 
33 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 17 5 7 8 16 13 14 15 12 22 
22 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 14 13 12 15 16 
16 1 2 3 9 9 4 5 6 7 8 9 10 10 19 17 10 
7 1 2 3 9 9 19 9 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
8 1 2 3 9 9 9 18 9 
30 1 2 3 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 11 10 13 15 14 12 16 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 18 9 
47 1 2 3 9 9 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 16 16 14 12 15 13 16 
39 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 5 17 7 8 10 5 17 7 8 10 10 11 10 17 5 7 8 16 14 12 13 15 22 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
7 1 2 20 3 20 18 9 
33 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 22 22 22 5 17 7 8 16 14 13 12 15 22 
3 1 2 18 
6 1 2 3 9 19 9 
4 1 2 18 20 
14 1 2 3 4 6 5 7 8 9 11 10 18 21 16 
26 1 2 3 9 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 14 15 12 13 22 
41 1 2 3 9 9 9 9 9 4 5 6 7 8 9 11 10 16 16 16 22 22 22 22 22 5 17 7 8 22 22 22 11 22 16 16 16 14 13 15 12 16 
25 1 2 3 20 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 14 13 15 12 16 
22 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
28 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 11 10 16 22 22 22 22 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
12 1 2 20 3 20 9 9 9 9 9 18 9 
4 1 2 18 20 
5 1 2 20 18 20 
3 1 2 18 
26 1 2 3 9 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 11 10 14 12 13 15 16 
3 1 2 18 
7 1 2 20 20 20 18 20 
3 1 2 18 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
36 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 16 17 5 7 8 22 22 22 11 22 16 14 13 12 15 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 16 14 13 12 15 16 
3 1 2 18 
24 1 2 3 20 4 9 9 9 9 9 9 9 9 9 5 6 7 8 9 10 10 17 19 10 
24 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 10 11 10 14 12 13 15 16 
24 1 2 3 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
7 1 2 20 3 20 18 9 
5 1 2 20 18 20 
17 1 2 3 9 9 9 4 5 6 7 8 9 10 10 17 19 10 
31 1 2 20 3 20 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 16 16 16 12 15 13 14 16 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
19 1 2 3 4 6 5 7 8 9 10 10 10 11 10 14 12 15 13 16 
6 1 2 3 20 18 9 
3 1 2 18 
33 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 16 17 5 7 8 22 22 22 22 11 22 16 13 14 15 12 16 
4 1 2 18 20 
21 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
7 1 2 3 9 9 18 9 
3 1 2 18 
3 1 2 18 
11 1 2 3 9 9 9 9 9 9 19 9 
10 1 2 3 20 9 9 9 9 19 9 
4 1 2 18 20 
3 1 2 18 
18 1 2 20 3 20 9 9 4 6 5 7 8 9 10 10 19 17 10 
37 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 16 16 16 16 16 18 21 16 
3 1 2 18 
19 1 2 3 9 4 6 5 7 8 9 10 11 10 16 12 15 14 13 16 
4 1 2 18 20 
16 1 2 3 4 6 5 7 8 9 11 10 14 15 12 13 16 
5 1 2 3 19 9 
4 1 2 18 20 
20 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 14 13 12 15 16 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 12 13 15 14 16 
7 1 2 3 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
28 1 2 3 4 5 6 7 8 9 10 10 10 5 17 7 8 10 17 5 7 8 10 10 10 10 17 19 10 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
19 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 17 19 10 
42 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 16 16 22 22 22 22 22 16 16 16 16 16 22 22 22 22 22 22 22 16 16 18 21 16 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
30 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 16 18 21 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 12 13 15 16 
7 1 2 3 20 4 18 9 
22 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 22 14 12 13 15 16 
3 1 2 18 
23 1 2 3 4 6 5 7 8 9 10 11 10 16 23 16 16 16 16 15 13 12 14 16 
8 1 2 3 20 9 9 19 9 
3 1 2 18 
20 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 11 10 21 18 16 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 18 9 
20 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 14 12 15 13 22 
4 1 2 18 20 
23 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 14 13 12 15 16 
6 1 2 3 20 18 9 
7 1 2 3 20 9 18 9 
3 1 2 18 
22 1 2 3 20 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 19 17 10 
17 1 2 3 9 9 4 5 6 7 8 9 10 11 10 21 18 16 
25 1 2 3 4 6 5 7 8 9 10 10 5 17 7 8 10 10 10 11 10 16 22 18 21 16 
4 1 2 18 20 
24 1 2 20 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 22 14 12 13 15 16 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 
37 1 2 3 20 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 18 21 22 
3 1 2 18 
23 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 14 15 13 12 16 
3 1 2 18 
4 1 2 18 20 
10 1 2 3 9 9 9 9 9 19 9 
4 1 2 18 20 
31 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 16 16 16 16 16 22 22 16 16 16 16 14 13 12 15 16 
3 1 2 18 
15 1 2 3 9 4 6 5 7 8 9 10 10 19 17 10 
30 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 11 10 16 22 22 22 16 16 14 12 13 15 16 
3 1 2 18 
5 1 2 3 19 9 
5 1 2 3 18 9 
36 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 16 5 17 7 8 16 11 22 13 14 12 15 16 
4 1 2 18 20 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
30 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 11 10 16 16 16 22 19 17 22 
3 1 2 18 
3 1 2 18 
18 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 17 19 10 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
31 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 17 5 7 8 22 22 11 22 14 13 15 12 16 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 14 15 13 12 16 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 19 9 
35 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 16 16 17 19 16 
3 1 2 18 
22 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 21 18 16 
3 1 2 18 
24 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 16 16 16 22 13 14 15 12 16 
3 1 2 18 
4 1 2 18 20 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
24 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
39 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 5 17 7 8 10 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
41 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 22 22 16 22 22 22 22 13 14 12 15 16 
3 1 2 18 
5 1 2 3 18 9 
25 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 16 18 21 16 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
25 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
21 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 19 17 10 
14 1 2 3 20 9 4 6 5 7 8 9 17 19 10 
5 1 2 3 18 9 
3 1 2 18 
24 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 11 10 16 16 14 12 15 13 16 
5 1 2 20 18 20 
34 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 11 10 16 22 22 22 22 17 5 7 8 16 12 13 15 14 22 
19 1 2 3 20 9 9 9 4 6 5 7 8 9 10 11 10 18 21 16 
4 1 2 18 20 
27 1 2 3 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 17 19 
3 1 2 18 
12 1 2 3 4 6 5 7 8 9 19 17 10 
3 1 2 18 
3 1 2 18 
5 1 2 23 18 23 
7 1 2 3 20 9 18 9 
35 1 2 3 4 5 6 7 8 9 10 10 10 11 10 5 17 7 8 16 22 22 22 22 22 22 22 22 22 11 22 14 12 13 15 16 
3 1 2 18 
15 1 2 3 9 4 5 6 7 8 9 10 10 17 19 10 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
12 1 2 20 3 20 9 9 9 9 9 18 9 
8 1 2 3 20 9 9 18 9 
9 1 2 3 20 9 9 9 9 19 
38 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 
36 1 2 3 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 22 15 13 14 12 16 
15 1 2 3 4 5 6 7 8 9 10 11 10 21 18 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
6 1 2 20 20 18 20 
4 1 2 18 20 
32 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 15 12 13 14 22 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 11 10 15 13 12 14 16 
18 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
15 1 2 3 4 6 5 7 8 9 10 11 10 21 18 16 
26 1 2 20 20 3 20 9 4 5 6 7 8 9 11 10 16 22 22 16 22 22 14 13 15 12 16 
21 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 14 15 13 12 16 
23 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 11 10 16 14 12 13 15 16 
17 1 2 3 4 5 6 7 8 9 10 10 10 11 10 21 18 16 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
7 1 2 20 20 20 18 20 
32 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 11 10 16 22 22 22 16 16 22 22 22 22 22 18 21 16 
19 1 2 20 3 20 9 9 4 5 6 7 8 9 11 10 16 21 18 22 
3 1 2 18 
23 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 14 15 13 12 16 
34 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 22 5 17 7 8 22 22 22 22 11 22 16 22 22 14 12 13 15 22 
48 1 2 20 3 20 9 4 6 5 7 8 9 17 5 7 8 10 5 17 7 8 10 5 17 7 8 10 10 10 10 11 10 16 16 22 22 22 22 17 5 7 8 16 14 12 15 13 22 
12 1 2 3 4 5 6 7 8 9 17 19 10 
7 1 2 3 9 4 19 9 
3 1 2 18 
5 1 2 20 18 20 
22 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 11 10 13 12 14 15 16 
32 1 2 3 9 9 9 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 11 10 16 22 22 22 16 22 19 17 22 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
10 1 2 20 20 3 20 9 9 18 9 
36 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
24 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
11 1 2 20 20 3 20 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
19 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 19 
32 1 2 20 20 3 20 4 5 6 7 8 9 11 10 16 16 22 22 17 5 7 8 22 22 22 22 22 14 13 15 12 22 
13 1 2 3 4 5 6 7 8 9 10 18 21 10 
23 1 2 3 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 17 19 10 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
15 1 2 3 4 6 5 7 8 9 10 11 10 21 18 16 
8 1 2 3 9 9 9 19 9 
24 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
26 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 22 21 18 22 
6 1 2 3 20 18 9 
14 1 2 3 9 4 6 5 7 8 9 10 17 19 10 
4 1 2 18 20 
6 1 2 3 20 18 9 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 13 14 12 15 16 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
4 1 2 18 20 
34 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 16 22 22 22 22 18 21 16 
36 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
9 1 2 20 3 20 9 9 18 9 
3 1 2 18 
12 1 2 3 4 6 5 7 8 9 19 17 10 
27 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
24 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
11 1 2 3 9 9 9 9 9 9 9 19 
30 1 2 3 4 6 5 7 8 9 10 10 17 5 7 8 10 10 10 10 11 10 16 16 16 22 15 13 12 14 22 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
27 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
24 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
20 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 14 13 15 12 16 
3 1 2 18 
25 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 14 12 13 15 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 19 9 
23 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 11 10 16 15 13 12 14 16 
3 1 2 18 
15 1 2 3 20 4 5 6 7 8 9 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 18 9 
30 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 16 22 16 15 12 14 13 16 
21 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 18 21 16 
53 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 21 18 16 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
23 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
6 1 2 20 20 18 20 
35 1 2 20 3 20 9 4 5 6 7 8 9 17 5 7 8 10 11 10 16 16 22 22 22 22 22 22 22 16 16 14 13 12 15 16 
6 1 2 3 9 19 9 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 10 10 17 19 10 
8 1 2 3 9 9 9 19 9 
65 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 16 16 16 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 5 17 7 8 16 17 5 7 8 22 22 22 22 22 11 22 16 15 13 14 12 16 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 20 19 9 
46 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 5 17 7 8 16 22 22 22 22 22 22 22 22 22 22 22 22 11 22 16 16 14 12 13 15 16 
37 1 2 20 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 5 17 7 8 10 5 17 7 8 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
21 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
11 1 2 3 9 9 9 9 9 9 9 19 
6 1 2 3 9 18 9 
3 1 2 18 
3 1 2 18 
24 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 16 16 16 14 15 13 12 16 
26 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 22 16 13 14 12 15 16 
10 1 2 3 20 9 9 9 9 18 9 
6 1 2 3 9 19 9 
5 1 2 3 19 9 
31 1 2 3 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 22 19 17 22 
5 1 2 3 19 9 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
14 1 2 3 20 9 9 9 9 9 9 9 9 19 9 
6 1 2 3 20 19 9 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 19 10 
36 1 2 3 4 9 6 5 7 8 9 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 14 13 15 12 16 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 19 17 10 
3 1 2 18 
9 1 2 3 9 9 9 9 9 19 
3 1 2 18 
4 1 2 18 20 
24 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 13 15 14 12 16 
18 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 21 18 16 
3 1 2 18 
17 1 2 3 20 4 6 5 7 8 9 10 10 10 10 17 19 10 
3 1 2 18 
7 1 2 3 20 9 18 9 
5 1 2 3 19 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 20 4 18 9 
23 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
20 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 11 10 21 18 16 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 11 10 16 16 21 18 16 
22 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 21 18 16 
4 1 2 18 20 
21 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
28 1 2 3 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 11 10 16 13 14 15 12 16 
36 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 16 16 22 22 22 22 22 22 17 5 7 8 22 22 11 22 14 12 13 15 16 
23 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 16 21 18 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 18 9 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 13 14 12 15 16 
6 1 2 3 20 18 9 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 21 18 16 
4 1 2 18 20 
22 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
8 1 2 3 9 9 9 19 9 
3 1 2 18 
28 1 2 3 4 5 6 7 8 9 10 10 11 10 16 17 5 7 8 16 22 22 11 22 14 15 13 12 16 
3 1 2 18 
35 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 16 16 21 18 16 
25 1 2 3 20 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 10 10 17 10 19 
4 1 2 18 20 
5 1 2 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
18 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 21 18 16 
3 1 2 18 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
5 1 2 3 18 9 
4 1 2 18 20 
4 1 2 18 20 
20 1 2 3 20 4 5 6 7 8 9 10 5 17 7 8 10 10 19 17 10 
30 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 16 17 5 7 8 16 14 12 13 15 22 
12 1 2 3 4 5 6 7 8 9 19 17 10 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
46 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 5 17 7 8 10 5 17 7 8 10 10 11 10 16 16 22 22 22 22 16 22 22 22 22 22 14 13 12 15 16 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
20 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 14 12 15 13 16 
15 1 2 3 9 4 5 6 7 8 9 10 10 17 19 10 
39 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 16 16 16 17 5 7 8 22 22 22 22 22 22 11 22 12 14 13 15 16 
40 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 17 5 7 8 10 10 5 17 7 8 10 10 10 10 10 10 10 17 5 7 8 10 10 11 10 
23 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 21 18 16 
16 1 2 3 4 5 6 7 8 9 11 10 14 12 15 13 16 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
17 1 2 3 9 4 5 6 7 8 9 10 11 10 16 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
21 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 12 14 13 15 16 
4 1 2 18 20 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
19 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
23 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
14 1 2 3 4 5 6 7 8 9 10 10 17 19 10 
17 1 2 3 9 9 9 4 5 6 7 8 9 10 10 17 19 10 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
24 1 2 3 4 5 6 7 8 9 5 17 7 8 10 11 10 16 16 16 12 13 15 14 16 
23 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 21 18 16 
17 1 2 3 9 9 9 9 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 18 9 
56 1 2 3 20 4 5 6 7 8 9 10 5 17 7 8 10 5 17 7 8 10 10 5 17 7 8 10 17 5 7 8 10 10 10 10 10 10 11 10 16 16 22 22 22 22 22 17 5 7 8 16 14 13 12 15 22 
9 1 2 20 20 20 20 20 18 20 
5 1 2 20 18 20 
30 1 2 20 3 20 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 16 13 14 15 12 16 
3 1 2 18 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 11 10 16 21 18 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
29 1 2 20 20 3 20 9 4 5 6 7 8 9 10 10 10 10 17 5 7 8 10 10 10 11 10 21 18 16 
19 1 2 20 3 20 4 5 6 7 8 9 10 11 10 14 15 13 12 16 
3 1 2 18 
4 1 2 18 20 
15 1 2 3 4 5 6 7 8 9 10 11 10 18 21 16 
5 1 2 20 18 20 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 15 13 12 16 
29 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 14 12 13 15 16 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
5 1 2 20 18 20 
24 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 17 19 10 
25 1 2 3 20 9 4 5 6 7 8 9 10 5 17 7 8 10 10 11 10 16 16 18 21 16 
5 1 2 3 18 9 
16 1 2 3 9 9 9 9 4 6 5 7 8 9 19 17 10 
3 1 2 18 
33 1 2 3 4 6 5 7 8 9 10 10 17 5 7 8 10 11 10 16 22 17 5 7 8 22 22 11 22 12 13 15 14 16 
18 1 2 3 20 4 6 5 7 8 9 10 11 10 13 14 12 15 16 
3 1 2 18 
10 1 2 3 20 9 9 9 9 18 9 
19 1 2 3 9 4 6 5 7 8 9 11 10 16 16 14 13 12 15 16 
12 1 2 3 4 5 6 7 8 9 17 19 10 
9 1 2 3 20 9 9 4 18 9 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
10 1 2 3 20 9 9 9 9 19 9 
4 1 2 18 20 
25 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 16 22 22 16 16 14 13 12 15 16 
6 1 2 3 9 18 9 
3 1 2 18 
19 1 2 20 3 20 9 4 6 5 7 8 9 10 10 11 10 21 18 16 
35 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 5 17 7 8 10 5 17 7 8 10 10 10 10 10 17 19 
4 1 2 18 20 
11 1 2 3 20 9 9 9 9 9 19 9 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 11 10 18 21 16 
6 1 2 3 9 18 9 
3 1 2 18 
13 1 2 20 20 20 20 20 3 20 9 9 18 9 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 13 12 14 15 16 
6 1 2 20 20 18 20 
7 1 2 3 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
21 1 2 20 3 20 9 4 6 5 7 8 9 10 10 11 10 14 12 15 13 16 
4 1 2 18 20 
6 1 2 20 20 18 20 
5 1 2 20 18 20 
28 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 14 12 13 15 16 
16 1 2 20 20 3 20 9 9 9 9 9 9 9 9 19 9 
5 1 2 20 18 20 
7 1 2 20 3 20 18 9 
22 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 21 18 16 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 19 9 
7 1 2 3 20 9 18 9 
19 1 2 20 3 20 4 6 5 7 8 9 10 11 10 15 13 12 14 16 
9 1 2 3 20 9 9 9 19 9 
3 1 2 18 
25 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 16 14 15 12 13 16 
8 1 2 3 9 9 9 9 19 
3 1 2 18 
35 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
22 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
23 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 
3 1 2 18 
23 1 2 20 20 20 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
27 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 16 22 22 22 22 16 16 12 13 14 15 16 
5 1 2 20 18 20 
4 1 2 18 20 
53 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 22 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 17 19 22 
42 1 2 20 20 20 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 16 17 5 7 8 22 22 22 22 22 22 11 22 14 15 13 12 16 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
23 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 16 21 18 16 
3 1 2 18 
32 1 2 3 20 9 4 6 5 7 8 9 10 10 11 10 16 23 23 23 16 22 22 22 22 22 22 16 14 12 13 15 16 
48 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 16 22 22 22 16 16 16 22 22 22 22 22 22 16 21 18 16 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
6 1 2 3 20 18 9 
4 1 2 18 20 
31 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 14 13 12 15 16 
4 1 2 18 20 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 18 21 16 
30 1 2 3 20 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
14 1 2 3 20 4 5 6 7 8 9 10 19 17 10 
4 1 2 18 20 
26 1 2 3 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 11 10 16 14 12 13 15 16 
8 1 2 3 20 9 9 18 9 
36 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
21 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 16 16 16 21 18 22 
17 1 2 3 20 4 6 5 7 8 9 10 11 10 16 21 18 16 
3 1 2 18 
3 1 2 18 
39 1 2 20 20 20 20 3 20 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 10 11 10 16 16 22 22 22 16 13 14 15 12 16 
5 1 2 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
20 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 14 12 15 13 16 
37 1 2 3 20 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 16 16 16 22 22 22 16 5 17 7 8 16 13 14 15 12 22 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
21 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 19 10 
5 1 2 3 18 9 
11 1 2 3 20 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 20 18 9 
14 1 2 3 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
21 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 14 15 13 12 16 
4 1 2 18 20 
5 1 2 3 19 9 
4 1 2 18 20 
19 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 19 17 10 
13 1 2 3 20 4 6 5 7 8 9 17 19 10 
33 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 16 22 22 22 22 22 22 16 16 22 22 22 14 15 12 13 16 
12 1 2 20 3 20 9 9 9 9 9 9 19 
38 1 2 20 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 14 13 15 12 16 
5 1 2 3 18 9 
4 1 2 18 20 
6 1 2 20 23 18 23 
3 1 2 18 
3 1 2 18 
21 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 16 14 13 12 15 16 
7 1 2 3 20 9 18 9 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
25 1 2 3 20 9 4 6 5 7 8 9 10 11 10 16 16 16 22 22 16 13 14 15 12 16 
4 1 2 18 20 
33 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 16 22 17 5 7 8 22 22 22 11 22 16 12 13 15 14 16 
4 1 2 18 20 
30 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 16 22 22 22 22 21 18 16 
4 1 2 18 20 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
16 1 2 3 20 9 9 9 4 6 5 7 8 9 19 17 10 
4 1 2 18 20 
19 1 2 3 20 4 5 6 7 8 9 10 11 10 16 16 16 17 19 22 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
42 1 2 3 9 4 6 5 7 8 9 10 10 10 5 17 7 8 10 10 5 17 7 8 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 10 
3 1 2 18 
5 1 2 20 18 20 
4 1 2 18 20 
19 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
19 1 2 3 20 4 6 5 7 8 9 5 17 7 8 10 10 19 17 10 
19 1 2 3 20 4 5 6 7 8 9 11 10 16 16 13 12 15 14 16 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
37 1 2 3 9 4 6 5 7 8 9 10 10 10 5 17 7 8 10 10 10 11 10 17 5 7 8 16 22 22 22 11 22 13 14 12 15 16 
13 1 2 3 20 9 9 9 9 9 9 9 9 19 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 10 19 17 
8 1 2 3 20 9 9 19 9 
20 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 13 14 12 15 16 
5 1 2 20 18 20 
26 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 16 14 12 13 15 16 
17 1 2 3 9 4 6 5 7 8 9 11 10 13 14 15 12 16 
21 1 2 20 20 3 20 4 5 6 7 8 9 10 10 11 10 15 12 14 13 16 
6 1 2 20 23 18 23 
3 1 2 18 
5 1 2 20 18 20 
8 1 2 20 3 20 9 19 9 
28 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 12 13 15 14 16 
4 1 2 18 20 
25 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 15 14 12 13 16 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 20 18 20 
26 1 2 20 3 20 9 4 5 6 7 8 9 10 10 11 10 16 16 22 16 22 13 12 14 15 16 
5 1 2 20 18 20 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 19 9 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
25 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 17 19 
11 1 2 3 20 9 9 9 9 9 19 9 
21 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 16 14 13 15 12 16 
30 1 2 3 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 14 13 12 15 16 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
8 1 2 3 20 9 9 18 9 
7 1 2 3 20 9 18 9 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
9 1 2 3 20 9 9 9 18 9 
4 1 2 18 20 
22 1 2 3 20 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
5 1 2 3 19 9 
19 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 19 17 10 
23 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 18 21 16 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
16 1 2 3 20 4 6 5 7 8 9 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
23 1 2 20 3 20 4 5 6 7 8 9 10 11 10 16 16 22 22 14 13 12 15 16 
22 1 2 20 3 20 4 5 6 7 8 9 17 5 7 8 10 10 11 10 21 18 16 
24 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 16 22 22 12 14 15 13 16 
15 1 2 3 4 5 6 7 8 9 10 10 10 19 17 10 
9 1 2 3 20 9 9 9 18 9 
12 1 2 20 3 20 9 9 9 9 9 9 19 
26 1 2 3 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 19 17 
3 1 2 18 
16 1 2 3 20 9 4 6 5 7 8 9 10 10 19 17 10 
5 1 2 20 18 20 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 14 13 12 15 16 
12 1 2 3 9 9 9 9 9 9 9 9 19 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 4 9 9 9 19 
4 1 2 18 20 
36 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 10 10 11 10 16 16 22 14 15 13 12 16 
22 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 21 18 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
9 1 2 3 20 9 9 9 18 9 
4 1 2 18 20 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
4 1 2 18 20 
38 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 11 10 16 22 22 22 17 5 7 8 16 14 13 12 15 22 
20 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 13 14 12 15 16 
21 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 17 19 10 
27 1 2 3 4 6 5 7 8 9 11 10 16 22 22 16 22 22 22 22 16 22 22 22 22 21 18 16 
33 1 2 3 20 4 6 5 7 8 9 10 17 5 7 8 10 17 5 7 8 10 5 17 7 8 10 10 10 11 10 18 21 16 
31 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 16 16 16 16 14 15 13 12 16 
36 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 22 16 16 22 22 22 5 17 7 8 22 22 22 11 22 14 12 13 15 16 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
15 1 2 3 4 5 6 7 8 9 10 10 10 10 19 17 
6 1 2 20 20 18 20 
4 1 2 18 20 
28 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 5 17 7 8 10 11 10 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 17 19 
63 1 2 3 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 17 5 7 8 10 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 17 19 22 
22 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
43 1 2 3 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 16 16 22 22 22 22 22 16 16 22 22 22 14 12 13 15 16 
28 1 2 3 20 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 11 10 21 18 16 
4 1 2 18 20 
22 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 22 22 14 13 12 15 16 
28 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 16 16 22 22 22 22 16 13 14 12 15 16 
8 1 2 3 9 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
6 1 2 20 20 18 20 
5 1 2 3 19 9 
4 1 2 18 20 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 12 13 14 15 16 
45 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 10 10 10 10 10 10 10 10 10 10 10 10 10 10 
14 1 2 3 4 5 6 7 8 9 10 10 17 19 10 
21 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 19 17 
14 1 2 3 20 4 5 6 7 8 9 10 21 18 10 
32 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 17 5 7 8 10 10 11 10 17 19 16 
16 1 2 3 4 5 6 7 8 9 10 10 11 10 19 17 16 
19 1 2 3 20 9 4 5 6 7 8 9 10 11 10 13 12 14 15 16 
4 1 2 18 20 
14 1 2 3 9 4 5 6 7 8 9 10 19 17 10 
21 1 2 3 20 4 5 6 7 8 9 11 10 16 16 22 16 12 14 13 15 16 
30 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 5 17 7 8 16 13 14 12 15 22 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
6 1 2 20 20 18 20 
7 1 2 3 20 4 19 9 
5 1 2 20 18 20 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
30 1 2 3 20 9 9 9 9 9 9 9 9 4 6 5 7 8 9 11 10 16 22 22 22 22 13 14 15 12 16 
12 1 2 20 3 20 9 9 9 9 9 9 19 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
5 1 2 3 18 9 
25 1 2 3 20 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
5 1 2 3 18 9 
7 1 2 3 20 4 18 9 
5 1 2 20 18 20 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
22 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
34 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 11 10 5 17 7 8 16 22 22 22 11 22 16 16 13 14 15 12 16 
6 1 2 3 20 18 9 
17 1 2 3 20 4 5 6 7 8 9 11 10 13 12 15 14 16 
23 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
21 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 16 15 13 12 14 16 
5 1 2 20 18 20 
3 1 2 18 
6 1 2 3 20 18 9 
22 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 18 21 16 
22 1 2 3 20 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 19 17 10 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
37 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 16 16 22 5 17 7 8 22 22 22 22 11 22 14 13 12 15 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
16 1 2 3 4 5 6 7 8 9 10 11 10 16 18 21 16 
41 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 5 17 7 8 10 11 10 16 16 22 22 22 16 16 22 22 22 22 22 17 19 22 
4 1 2 18 20 
59 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 11 22 16 22 22 16 16 16 14 13 12 15 16 
4 1 2 18 20 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 19 9 
7 1 2 3 9 9 19 9 
3 1 2 18 
33 1 2 20 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 16 5 17 7 8 16 14 13 12 15 22 
3 1 2 18 
3 1 2 18 
19 1 2 3 9 4 5 6 7 8 9 10 11 10 16 14 15 12 13 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
31 1 2 3 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 11 10 13 12 15 14 16 
4 1 2 18 20 
24 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 13 14 12 15 16 
4 1 2 18 20 
24 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 19 17 10 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
31 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 11 10 16 16 16 13 14 15 12 16 
8 1 2 3 9 9 9 19 9 
32 1 2 3 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 11 10 21 18 16 
5 1 2 3 18 9 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 15 14 12 13 16 
27 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 10 11 10 16 16 16 14 13 15 12 16 
3 1 2 18 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
17 1 2 3 4 6 5 7 8 9 10 10 11 10 16 21 18 16 
3 1 2 18 
22 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 18 21 16 
5 1 2 3 18 9 
37 1 2 3 9 4 6 5 7 8 9 10 10 10 17 5 7 8 10 10 10 11 10 16 16 16 22 22 22 22 16 16 16 14 12 13 15 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 16 23 21 18 16 
21 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 14 12 13 15 16 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 21 18 16 
4 1 2 18 20 
6 1 2 20 20 18 20 
3 1 2 18 
4 1 2 18 20 
26 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 21 18 16 
29 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 17 19 10 
4 1 2 18 20 
29 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 11 10 18 21 16 
17 1 2 3 4 5 6 7 8 9 10 11 10 12 14 13 15 16 
25 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 10 19 17 10 
35 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 16 16 16 22 22 16 16 16 16 16 16 14 12 13 15 16 
39 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 16 22 22 22 16 17 5 7 8 16 15 13 12 14 22 
3 1 2 18 
6 1 2 3 20 18 9 
24 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
24 1 2 20 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 21 18 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 15 13 12 14 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
25 1 2 3 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 11 10 21 18 16 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
17 1 2 3 20 9 9 4 5 6 7 8 9 10 10 19 17 10 
6 1 2 3 9 19 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
4 1 2 18 20 
26 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 14 15 12 13 16 
33 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 11 10 18 21 16 
4 1 2 18 20 
25 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 21 18 16 
28 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
4 1 2 18 20 
53 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
4 1 2 18 20 
26 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 16 14 12 15 13 16 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 10 
20 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 15 13 12 14 16 
28 1 2 3 20 4 6 5 7 8 9 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 19 17 
20 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 10 19 17 10 
22 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 16 22 14 13 15 12 16 
26 1 2 20 3 20 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 19 17 10 
11 1 2 20 20 20 3 20 9 9 19 9 
6 1 2 3 9 18 9 
45 1 2 3 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 11 10 16 16 22 22 22 22 16 16 17 5 7 8 16 22 22 22 11 22 16 14 13 12 15 16 
16 1 2 3 4 5 6 7 8 9 11 10 12 13 15 14 16 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 10 17 19 
22 1 2 3 4 5 6 7 8 9 11 10 16 16 16 22 22 22 14 13 15 12 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
7 1 2 20 3 20 18 9 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
21 1 2 3 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 17 19 10 
5 1 2 20 18 20 
33 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
11 1 2 3 9 9 9 9 4 9 19 9 
5 1 2 3 18 9 
5 1 2 3 19 9 
36 1 2 20 3 20 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 16 16 16 16 13 14 12 15 16 
5 1 2 3 19 9 
3 1 2 18 
5 1 2 3 19 9 
5 1 2 3 18 9 
5 1 2 3 19 9 
5 1 2 20 18 20 
5 1 2 3 19 9 
5 1 2 3 19 9 
5 1 2 3 19 9 
5 1 2 3 19 9 
5 1 2 3 19 9 
7 1 2 3 20 9 18 9 
5 1 2 3 19 9 
4 1 2 18 20 
6 1 2 3 20 18 9 
6 1 2 3 20 18 9 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
20 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 21 18 22 
5 1 2 3 18 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 17 19 22 
4 1 2 18 20 
22 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 10 
16 1 2 3 4 6 5 7 8 9 11 10 15 12 14 13 16 
4 1 2 18 20 
48 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 17 5 7 8 10 10 10 10 10 11 10 17 5 7 8 16 11 22 16 16 22 22 22 22 22 16 22 22 12 13 15 14 16 
51 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 17 5 7 8 22 22 22 11 22 16 16 22 22 22 22 22 22 22 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
43 1 2 3 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 10 11 10 16 16 16 16 16 16 16 22 22 22 22 22 22 22 16 16 13 12 14 15 16 
11 1 2 3 9 9 9 9 9 9 9 19 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 17 19 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
15 1 2 3 9 4 6 5 7 8 9 10 10 19 17 10 
18 1 2 3 20 4 5 6 7 8 9 10 11 10 14 15 13 12 16 
7 1 2 3 20 9 18 9 
30 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
27 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 17 19 
26 1 2 3 20 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 14 12 13 15 16 
6 1 2 3 20 18 9 
21 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
7 1 2 20 20 20 18 20 
30 1 2 20 20 20 20 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 11 10 12 13 15 14 16 
25 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 16 16 22 22 16 14 12 13 15 16 
3 1 2 18 
24 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 16 14 13 15 12 16 
3 1 2 18 
21 1 2 20 20 3 20 9 9 9 9 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
22 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 11 10 14 13 12 15 16 
25 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 11 10 18 21 16 
45 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 16 16 16 16 22 22 22 16 16 16 16 22 22 22 16 5 17 7 8 16 14 12 13 15 22 
9 1 2 3 20 9 9 9 18 9 
22 1 2 3 20 4 6 5 7 8 9 10 10 11 10 14 12 13 15 16 16 16 16 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
4 1 2 18 20 
18 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 20 9 4 6 5 7 8 9 10 11 10 16 16 21 18 16 
4 1 2 18 20 
14 1 2 3 4 6 5 7 8 9 10 10 17 19 10 
4 1 2 18 20 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
7 1 2 3 20 9 19 9 
6 1 2 3 20 19 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 18 9 
6 1 2 3 20 18 9 
3 1 2 18 
7 1 2 3 20 9 19 9 
68 1 2 3 20 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 11 10 16 16 22 22 22 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 5 17 7 8 22 22 14 13 12 15 22 
26 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 16 16 22 22 22 15 13 12 14 16 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
20 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 13 15 14 12 16 
4 1 2 18 20 
31 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 5 17 7 8 10 10 10 11 10 16 22 22 22 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
3 1 2 18 
18 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 18 21 16 
3 1 2 18 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
72 1 2 3 20 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 16 22 22 22 17 5 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 16 16 14 15 13 12 16 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
3 1 2 18 
4 1 2 18 20 
5 1 2 3 18 9 
32 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 5 17 7 8 10 10 10 11 10 14 15 13 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
8 1 2 3 9 9 9 9 19 
19 1 2 3 20 4 5 6 7 8 9 10 10 11 10 14 13 15 12 16 
3 1 2 18 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 16 15 14 12 13 16 
4 1 2 18 20 
5 1 2 20 18 20 
38 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 13 14 15 12 16 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 17 19 10 
22 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 10 
7 1 2 3 20 4 19 9 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
24 1 2 3 4 6 5 7 8 9 10 10 10 10 10 5 17 7 8 10 10 10 10 11 10 
25 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
31 1 2 3 4 5 6 7 8 9 5 17 7 8 10 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 19 17 
18 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 18 21 16 
8 1 2 3 9 9 9 9 19 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
34 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 5 17 7 8 22 22 22 22 22 22 22 11 22 13 12 14 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
26 1 2 3 20 9 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 10 17 19 10 
13 1 2 3 9 4 6 5 7 8 9 19 17 10 
14 1 2 3 20 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
9 1 2 23 23 20 20 23 18 20 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
5 1 2 23 18 23 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
26 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
29 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
21 1 2 3 9 9 4 5 6 7 8 9 11 10 16 16 16 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 4 5 6 7 8 9 11 10 16 23 16 22 22 15 14 12 13 16 
21 1 2 3 4 6 5 7 8 9 10 10 10 5 17 7 8 10 10 10 10 10 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 15 13 12 16 
9 1 2 20 20 3 20 9 18 9 
16 1 2 3 9 9 9 9 4 5 6 7 8 9 19 17 10 
10 1 2 3 9 9 9 9 9 19 9 
28 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 16 16 16 16 13 14 12 15 16 
27 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 13 14 12 15 16 
21 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
33 1 2 20 3 20 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 16 16 5 17 7 8 16 14 12 15 13 22 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
10 1 2 3 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
26 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 16 16 14 12 13 15 16 
5 1 2 20 18 20 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
7 1 2 3 20 9 18 9 
21 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 16 14 13 15 12 16 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 14 12 13 15 16 
19 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
26 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 14 12 13 15 16 
26 1 2 3 9 4 5 6 7 8 9 10 10 10 10 17 5 7 8 10 11 10 13 15 12 14 16 
16 1 2 3 20 4 6 5 7 8 9 10 10 10 17 19 10 
3 1 2 18 
10 1 2 20 3 20 9 9 9 18 9 
7 1 2 3 20 9 18 9 
18 1 2 20 20 20 20 20 3 20 4 5 6 7 8 9 17 19 10 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
3 1 2 18 
36 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 11 10 16 16 16 16 16 16 22 22 22 22 14 12 15 13 16 
3 1 2 18 
30 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 11 10 17 5 7 8 16 12 14 13 15 22 
17 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 19 17 
3 1 2 18 
31 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 16 16 21 18 16 
21 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 19 17 22 
4 1 2 18 20 
20 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 17 19 10 
7 1 2 3 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
7 1 2 3 20 9 18 9 
5 1 2 20 18 20 
17 1 2 3 9 4 5 6 7 8 9 10 11 10 16 18 21 16 
4 1 2 18 20 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
38 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 16 16 16 22 22 5 17 7 8 22 22 22 22 22 11 22 16 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
24 1 2 3 20 9 4 5 6 7 8 9 11 10 16 16 22 22 22 22 15 13 12 14 16 
4 1 2 18 20 
30 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 13 14 15 12 16 
13 1 2 3 9 4 5 6 7 8 9 17 19 10 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
20 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 13 14 12 15 16 
7 1 2 3 20 9 18 9 
17 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 17 19 
58 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 11 22 16 12 13 15 14 16 
26 1 2 3 20 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 11 10 21 18 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
28 1 2 3 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 10 10 10 11 10 14 15 12 13 16 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
7 1 2 3 9 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 9 18 9 
5 1 2 20 18 20 
26 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 16 16 14 12 13 15 16 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
31 1 2 3 4 6 5 7 8 9 17 5 7 8 10 11 10 16 22 22 22 22 22 16 22 22 16 14 12 13 15 16 
8 1 2 3 9 9 9 18 9 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
15 1 2 3 20 9 4 6 5 7 8 9 10 10 19 17 
6 1 2 3 9 19 9 
24 1 2 3 9 9 9 4 6 5 7 8 9 11 10 16 16 16 16 22 22 22 21 18 16 
9 1 2 3 9 9 9 9 19 9 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 16 14 13 15 12 16 
21 1 2 3 9 9 9 4 6 5 7 8 9 10 10 11 10 14 12 13 15 16 
3 1 2 18 
20 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 19 17 
5 1 2 3 18 9 
21 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 13 12 14 15 16 
4 1 2 18 20 
26 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 11 10 13 12 14 15 16 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 14 12 15 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
24 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 17 19 10 
28 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 16 16 16 16 22 22 22 16 13 14 15 12 16 
4 1 2 18 20 
3 1 2 18 
9 1 2 3 9 9 9 4 19 9 
27 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
23 1 2 3 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 21 18 16 
6 1 2 3 20 19 9 
4 1 2 18 20 
32 1 2 3 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
6 1 2 3 9 19 9 
20 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 14 12 13 15 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 20 9 18 9 
34 1 2 3 20 9 4 6 5 7 8 9 10 10 10 5 17 7 8 10 10 11 10 16 22 22 22 22 22 22 22 22 18 21 22 
4 1 2 18 20 
25 1 2 3 9 9 9 9 9 4 5 6 7 8 9 11 10 16 22 22 22 14 12 15 13 16 
3 1 2 18 
3 1 2 18 
29 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
15 1 2 3 9 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
28 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 14 15 13 12 22 
43 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 5 17 7 8 10 11 10 16 16 22 22 22 16 22 22 22 22 22 22 22 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
20 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 14 15 12 13 16 
8 1 2 3 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
24 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 16 22 22 13 12 14 15 22 
6 1 2 3 20 19 9 
11 1 2 3 20 9 9 9 9 9 18 9 
13 1 2 3 9 4 6 5 7 8 9 17 19 10 
3 1 2 18 
27 1 2 3 20 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 9 9 9 19 
7 1 2 3 9 9 18 9 
17 1 2 3 20 4 6 5 7 8 9 10 10 11 10 18 21 16 
9 1 2 3 9 9 9 9 9 19 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
5 1 2 3 18 9 
4 1 2 18 20 
13 1 2 3 9 4 5 6 7 8 9 17 19 10 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
37 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 17 5 7 8 10 10 11 10 16 22 22 15 14 13 12 16 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
13 1 2 3 9 4 6 5 7 8 9 17 19 10 
4 1 2 18 20 
4 1 2 18 20 
25 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 16 22 22 16 22 13 14 15 12 16 
40 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 5 17 7 8 22 22 22 22 22 22 22 11 22 13 14 12 15 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
22 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 16 22 22 22 18 21 16 
8 1 2 3 9 9 9 9 19 
25 1 2 3 9 9 4 6 5 7 8 9 10 5 17 7 8 10 10 11 10 13 14 15 12 16 
21 1 2 20 3 20 9 9 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
19 1 2 3 9 4 6 5 7 8 9 10 10 11 10 14 13 12 15 16 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 12 15 13 16 
3 1 2 18 
35 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 21 18 16 
52 1 2 20 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 19 17 16 
31 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 17 5 7 8 10 11 10 16 16 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
6 1 2 20 20 18 20 
3 1 2 18 
23 1 2 3 4 6 5 7 8 9 10 11 10 16 16 16 22 22 22 14 12 15 13 16 
3 1 2 18 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
11 1 2 3 9 9 9 9 9 9 18 9 
20 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 21 18 22 
4 1 2 18 20 
33 1 2 3 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 5 17 7 8 16 14 12 13 15 22 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
19 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
34 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 16 22 22 16 22 22 22 22 22 22 16 14 13 15 12 16 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 13 14 12 15 16 
33 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 16 16 22 22 22 13 14 12 15 16 
15 1 2 20 20 20 20 20 20 20 20 20 3 20 18 9 
4 1 2 18 20 
7 1 2 20 3 20 18 9 
6 1 2 20 20 18 20 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 19 17 
31 1 2 3 4 5 6 7 8 9 11 10 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 14 12 13 15 22 
18 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 17 19 10 
8 1 2 20 20 3 20 18 9 
19 1 2 3 4 5 6 7 8 9 5 17 7 8 10 11 10 21 18 16 
4 1 2 18 20 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
4 1 2 18 20 
17 1 2 3 4 6 5 7 8 9 11 10 16 14 13 15 12 16 
37 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 11 10 5 17 7 8 16 22 11 22 16 22 22 22 22 22 13 12 14 15 16 
5 1 2 3 19 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 19 9 
30 1 2 3 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 11 10 16 22 15 13 14 12 16 
3 1 2 18 
46 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 5 17 7 8 10 17 5 7 8 10 10 17 5 7 8 10 10 10 10 11 10 16 23 16 16 22 21 18 22 
22 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
5 1 2 20 18 20 
24 1 2 3 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 21 18 16 
3 1 2 18 
3 1 2 18 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
43 1 2 20 20 3 20 9 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 11 10 16 22 22 22 16 22 22 22 22 22 22 22 22 15 13 12 14 16 
25 1 2 3 4 6 5 7 8 9 5 17 7 8 10 17 5 7 8 10 10 10 10 17 19 10 
30 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 11 10 5 17 7 8 16 14 13 15 12 22 
16 1 2 3 4 5 6 7 8 9 10 10 11 10 19 17 16 
25 1 2 3 4 9 9 9 9 5 6 7 8 9 10 10 10 10 11 10 16 13 14 15 12 16 
6 1 2 20 20 18 20 
3 1 2 18 
8 1 2 20 3 20 9 18 9 
23 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 18 21 16 
8 1 2 20 3 20 9 18 9 
6 1 2 23 23 18 23 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 14 13 15 12 16 
17 1 2 3 4 6 5 7 8 9 10 10 10 11 10 21 18 16 
23 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
34 1 2 3 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 21 18 22 
20 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 15 14 12 13 16 
43 1 2 3 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 16 16 16 22 22 22 16 16 16 16 16 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
9 1 2 3 20 9 9 9 9 19 
22 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 11 10 21 18 16 
40 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 16 16 16 16 16 5 17 7 8 22 22 22 22 22 22 22 22 11 22 13 12 14 15 16 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
8 1 2 3 20 9 9 18 9 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 11 10 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
8 1 2 3 9 9 9 9 19 
28 1 2 3 20 9 4 5 6 7 8 9 10 10 10 11 10 16 16 17 5 7 8 16 14 12 13 15 22 
6 1 2 3 20 18 9 
13 1 2 3 9 4 6 5 7 8 9 17 19 10 
38 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 10 
8 1 2 3 9 9 9 18 9 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 14 12 15 16 
30 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 11 10 16 22 18 21 22 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 13 14 12 15 16 
4 1 2 18 20 
29 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 
29 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 11 10 16 22 22 16 22 22 14 13 15 12 16 
4 1 2 18 20 
9 1 2 3 20 9 9 9 9 19 
3 1 2 18 
7 1 2 3 20 9 19 9 
36 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 5 17 7 8 10 17 5 7 8 10 10 10 11 10 15 13 14 12 16 
3 1 2 18 
30 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 19 17 22 
3 1 2 18 
22 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 22 13 14 12 15 16 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
22 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 16 14 12 15 13 16 
24 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 12 14 13 15 16 
22 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 11 10 13 14 15 12 16 
12 1 2 3 20 9 9 9 9 9 9 9 19 
25 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 16 14 12 13 15 16 
18 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 17 19 10 
27 1 2 20 3 20 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 22 21 18 16 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 13 15 12 16 
43 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 17 5 7 8 10 10 17 5 7 8 10 10 10 10 17 5 7 8 10 10 10 10 
4 1 2 18 20 
19 1 2 3 20 9 4 6 5 7 8 9 10 10 10 11 10 21 18 16 
7 1 2 3 20 9 18 9 
18 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 19 17 22 
4 1 2 18 20 
4 1 2 18 20 
30 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 11 10 16 12 13 14 15 16 
24 1 2 20 20 20 20 3 20 9 4 5 6 7 8 9 10 10 11 10 15 14 12 13 16 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 14 15 13 12 16 
16 1 2 3 4 6 5 7 8 9 11 10 14 12 13 15 16 
24 1 2 3 20 9 4 6 5 7 8 9 10 11 10 16 16 22 22 22 22 16 19 17 16 
28 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 14 13 15 12 16 
29 1 2 3 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
36 1 2 3 20 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 14 12 13 15 16 
21 1 2 3 20 9 4 6 5 7 8 9 10 10 11 10 16 14 15 12 13 16 
4 1 2 18 20 
34 1 2 3 4 5 6 7 8 9 11 10 16 22 22 5 17 7 8 22 22 22 22 11 22 16 22 22 22 22 14 13 15 12 16 
37 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 22 22 22 22 22 16 22 22 16 16 22 16 16 16 16 16 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 18 9 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 3 19 9 
3 1 2 18 
11 1 2 20 20 3 20 9 9 9 19 9 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 13 14 12 15 16 
35 1 2 20 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 11 10 21 18 16 
29 1 2 3 4 6 5 7 8 9 11 10 17 5 7 8 16 22 22 22 22 22 11 22 16 14 12 15 13 16 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 14 12 13 15 22 
8 1 2 3 9 9 9 19 9 
25 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 5 17 7 8 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
9 1 2 20 20 20 20 20 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
24 1 2 3 9 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
21 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 16 12 14 15 13 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 19 17 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
6 1 2 20 20 18 20 
16 1 2 3 20 4 6 5 7 8 9 10 10 10 17 19 10 
19 1 2 3 4 6 5 7 8 9 11 10 16 22 22 14 13 12 15 16 
3 1 2 18 
39 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 11 10 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
27 1 2 20 3 20 9 9 4 6 5 7 8 9 10 11 10 16 16 16 22 22 22 13 12 15 14 16 
26 1 2 3 20 9 9 4 6 5 7 8 9 10 10 5 17 7 8 10 10 10 11 10 18 21 16 
15 1 2 3 4 5 6 7 8 9 10 11 10 18 21 16 
16 1 2 3 20 4 5 6 7 8 9 10 10 10 17 19 10 
19 1 2 3 20 9 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
23 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
12 1 2 3 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
39 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 5 17 7 8 10 10 10 11 10 16 16 22 22 5 17 7 8 22 14 12 13 15 22 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
27 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 22 22 22 13 15 12 14 16 
16 1 2 3 4 6 5 7 8 9 11 10 13 14 15 12 16 
6 1 2 3 20 18 9 
3 1 2 18 
39 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 11 10 16 22 22 22 12 14 13 15 16 
4 1 2 18 20 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 13 14 15 12 16 
35 1 2 3 20 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 16 22 22 22 16 22 22 22 14 13 15 12 16 
7 1 2 3 20 9 18 9 
23 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 11 10 13 14 12 15 16 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 21 18 16 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 3 9 4 9 6 5 7 8 9 10 10 10 10 10 10 10 17 19 
24 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 16 16 16 16 13 14 15 12 16 
11 1 2 3 9 9 9 9 9 9 9 19 
4 1 2 18 20 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
19 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 17 19 10 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
18 1 2 20 3 20 4 6 5 7 8 9 10 10 10 10 19 17 10 
30 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
7 1 2 3 20 9 19 9 
23 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 19 
23 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
35 1 2 3 20 9 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 22 22 22 22 17 5 7 8 16 14 13 12 15 22 
32 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 16 16 16 16 16 16 16 16 16 16 16 16 13 14 12 15 16 
3 1 2 18 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 17 19 10 
3 1 2 18 
14 1 2 3 9 9 4 6 5 7 8 9 19 17 10 
6 1 2 3 20 18 9 
22 1 2 3 4 6 5 7 8 9 10 10 10 10 10 11 10 16 12 15 14 13 16 
22 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 16 14 12 13 15 16 
4 1 2 18 20 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
23 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 15 14 13 12 16 
26 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 15 13 12 14 16 
26 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
24 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
31 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 16 16 22 22 22 22 22 14 15 13 12 16 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
24 1 2 3 4 6 5 7 8 9 10 10 17 5 7 8 10 10 11 10 13 12 14 15 16 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 11 10 21 18 16 
5 1 2 3 18 9 
18 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 18 21 16 
27 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 
16 1 2 3 4 6 5 7 8 9 11 10 14 13 12 15 16 
17 1 2 3 4 5 6 7 8 9 17 5 7 8 10 18 21 10 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 14 12 13 15 16 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
24 1 2 20 20 20 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
22 1 2 3 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 16 21 18 16 
3 1 2 18 
6 1 2 3 20 19 9 
36 1 2 20 20 3 20 9 4 6 5 7 8 9 10 10 11 10 16 16 22 5 17 7 8 22 22 22 22 22 22 22 11 22 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 16 21 18 16 
13 1 2 20 3 20 9 9 9 9 9 9 18 9 
8 1 2 20 20 20 20 18 20 
4 1 2 18 20 
16 1 2 3 20 9 9 4 6 5 7 8 9 10 19 17 10 
34 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 16 16 18 21 16 
43 1 2 3 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 5 17 7 8 10 10 17 5 7 8 10 10 10 11 10 16 16 22 22 22 13 14 15 12 16 
7 1 2 3 20 9 19 9 
19 1 2 3 20 9 4 5 6 7 8 9 10 10 10 11 10 21 18 16 
6 1 2 3 9 19 9 
3 1 2 18 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
3 1 2 18 
3 1 2 18 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
18 1 2 3 20 4 5 6 7 8 9 10 11 10 13 12 14 15 16 
22 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 17 19 
3 1 2 18 
17 1 2 3 20 4 5 6 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
24 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
6 1 2 3 20 18 9 
45 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 5 17 7 8 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 17 19 22 
3 1 2 18 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
24 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 16 14 15 13 12 16 
26 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
28 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 14 15 12 13 16 
9 1 2 3 9 9 9 9 19 9 
21 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
20 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 14 13 12 15 16 
25 1 2 3 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 11 10 13 14 12 15 16 
4 1 2 18 20 
11 1 2 3 20 9 9 9 9 9 18 9 
4 1 2 18 20 
21 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 10 10 10 17 19 10 
19 1 2 3 20 9 9 9 4 5 6 7 8 9 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
10 1 2 3 20 9 9 9 9 18 9 
5 1 2 20 18 20 
19 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 17 19 
32 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 17 5 7 8 22 22 22 11 22 21 18 16 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 4 6 5 7 8 9 10 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
30 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 
22 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 17 19 10 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 15 13 12 14 16 
19 1 2 3 4 6 5 7 8 9 10 10 10 11 10 15 13 12 14 16 
3 1 2 18 
5 1 2 3 19 9 
19 1 2 3 4 6 5 7 8 9 11 10 16 22 22 14 15 13 12 16 
3 1 2 18 
26 1 2 20 20 3 20 4 5 6 7 8 9 17 5 7 8 10 11 10 16 23 16 16 21 18 16 
28 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 11 10 16 5 17 7 8 16 15 14 12 13 22 
14 1 2 3 20 4 5 6 7 8 9 10 19 17 10 
4 1 2 18 20 
6 1 2 3 20 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
31 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 5 17 7 8 10 10 11 10 13 14 15 12 16 
4 1 2 18 20 
3 1 2 18 
5 1 2 20 18 20 
32 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 5 7 8 10 5 17 7 8 10 17 5 7 8 10 18 21 10 
51 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 22 22 22 22 22 22 22 22 18 21 16 
20 1 2 3 9 9 4 6 5 7 8 9 11 10 16 16 14 12 15 13 16 
3 1 2 18 
3 1 2 18 
8 1 2 20 3 20 9 18 9 
3 1 2 18 
28 1 2 3 20 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 17 19 10 
6 1 2 3 9 19 9 
7 1 2 3 20 9 18 9 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
5 1 2 23 18 23 
3 1 2 18 
3 1 2 18 
32 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 16 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
6 1 2 20 20 18 20 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
3 1 2 18 
16 1 2 3 9 9 4 6 5 7 8 9 10 10 19 17 10 
7 1 2 3 9 9 9 19 
39 1 2 3 20 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 16 16 16 16 16 16 16 22 22 22 22 22 22 22 22 14 12 15 13 16 
6 1 2 3 20 18 9 
3 1 2 18 
33 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 16 16 5 17 7 8 16 22 22 22 22 21 18 22 
23 1 2 3 20 4 6 5 7 8 9 11 10 16 16 16 22 22 16 12 14 13 15 16 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 14 12 15 13 16 
28 1 2 20 3 20 4 5 6 7 8 9 17 5 7 8 10 11 10 17 5 7 8 16 14 13 12 15 22 
3 1 2 18 
33 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 12 14 13 15 16 
5 1 2 3 18 9 
30 1 2 20 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 11 10 16 14 15 13 12 16 
7 1 2 3 20 9 18 9 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
6 1 2 20 20 18 20 
21 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 19 17 
14 1 2 20 20 3 20 9 9 9 9 9 9 9 19 
22 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
12 1 2 3 20 9 9 9 9 9 9 18 9 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
11 1 2 20 3 20 9 9 9 9 19 9 
29 1 2 3 20 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
20 1 2 3 4 6 5 7 8 9 11 10 16 16 16 22 22 22 18 21 16 
31 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 16 16 22 22 22 16 16 12 13 15 14 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
10 1 2 3 9 9 9 9 9 19 9 
20 1 2 3 4 5 6 7 8 9 11 10 16 22 22 16 22 16 21 18 16 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
7 1 2 3 20 9 18 9 
3 1 2 18 
24 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 14 13 12 15 16 
8 1 2 3 20 9 9 19 9 
19 1 2 3 9 9 9 9 4 5 6 7 8 9 11 10 16 21 18 16 
22 1 2 3 20 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 19 17 10 
24 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 18 21 16 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
43 1 2 3 20 4 5 6 7 8 9 10 10 11 10 5 17 7 8 16 22 22 11 22 16 22 22 5 17 7 8 22 22 17 5 7 8 22 22 14 12 13 15 22 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 9 4 5 6 7 8 9 11 10 14 13 12 15 16 
5 1 2 20 18 20 
5 1 2 3 19 9 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 19 17 
20 1 2 3 9 9 9 9 4 6 5 7 8 9 10 11 10 16 18 21 16 
20 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 11 10 18 21 16 
48 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 17 5 7 8 22 22 22 22 22 22 22 22 11 22 16 22 22 22 22 22 22 13 14 15 12 22 
10 1 2 3 9 9 9 9 9 19 9 
15 1 2 3 4 5 6 7 8 9 10 11 10 21 18 16 
17 1 2 3 9 9 9 9 4 6 5 7 8 9 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
42 1 2 20 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 17 5 7 8 10 17 5 7 8 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 
15 1 2 3 9 4 6 5 7 8 9 10 10 19 17 10 
4 1 2 18 20 
10 1 2 3 20 9 9 9 9 18 9 
5 1 2 3 19 9 
5 1 2 3 18 9 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
8 1 2 3 20 9 9 19 9 
17 1 2 3 4 5 6 7 8 9 10 11 10 13 15 12 14 16 
23 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
9 1 2 3 9 9 9 9 9 19 
3 1 2 18 
21 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 16 14 13 12 15 16 
19 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 17 19 10 
14 1 2 3 20 9 9 9 9 9 9 9 4 18 9 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 18 9 
14 1 2 3 9 9 4 5 6 7 8 9 19 17 10 
4 1 2 18 20 
3 1 2 18 
25 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 14 12 15 13 16 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
21 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
22 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
6 1 2 3 20 18 9 
6 1 2 3 20 19 9 
24 1 2 20 20 20 20 20 20 3 20 4 6 5 7 8 9 10 11 10 15 13 14 12 16 
37 1 2 3 4 9 9 9 9 9 9 9 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 17 5 7 8 10 10 11 10 18 21 16 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
31 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 10 10 10 11 10 14 13 12 15 16 
30 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 22 22 16 22 16 22 14 12 15 13 16 
5 1 2 3 18 9 
4 1 2 18 20 
16 1 2 3 20 9 4 5 6 7 8 9 11 10 21 18 16 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 13 14 12 15 16 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 18 9 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 19 17 
8 1 2 3 20 9 9 19 9 
4 1 2 18 20 
12 1 2 3 9 9 9 9 9 9 9 19 9 
14 1 2 3 20 9 9 9 9 9 9 9 9 18 9 
32 1 2 3 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 17 5 7 8 16 13 14 15 12 22 
4 1 2 18 20 
10 1 2 3 20 9 9 9 9 18 9 
4 1 2 18 20 
16 1 2 3 20 9 4 6 5 7 8 9 10 10 17 19 10 
3 1 2 18 
22 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 14 15 13 12 16 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
11 1 2 3 9 9 9 9 9 9 9 19 
4 1 2 18 20 
32 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 5 17 7 8 16 22 11 22 14 15 13 12 16 
3 1 2 18 
29 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 14 13 12 15 16 
31 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 16 23 16 16 22 22 22 22 16 16 16 14 12 15 13 16 
6 1 2 3 9 18 9 
22 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
15 1 2 3 20 9 4 5 6 7 8 9 10 19 17 10 
16 1 2 3 20 9 4 6 5 7 8 9 10 10 17 19 10 
15 1 2 3 20 9 4 6 5 7 8 9 10 17 19 10 
4 1 2 18 20 
30 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 12 13 15 14 16 
5 1 2 23 18 23 
3 1 2 18 
18 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 17 19 10 
19 1 2 3 20 9 4 6 5 7 8 9 10 11 10 13 14 15 12 16 
4 1 2 18 20 
34 1 2 3 20 9 9 4 6 5 7 8 9 10 10 17 5 7 8 10 10 10 10 11 10 16 22 22 16 16 12 14 13 15 16 
60 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 22 22 22 22 22 16 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 21 18 22 
6 1 2 3 4 19 9 
29 1 2 3 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 12 13 14 15 16 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
21 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
8 1 2 3 20 9 9 19 9 
46 1 2 3 9 9 9 9 9 4 9 5 6 7 8 9 5 17 7 8 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 16 22 22 16 16 22 22 22 22 21 18 16 
3 1 2 18 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
65 1 2 3 20 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 5 17 7 8 10 5 17 7 8 10 10 10 10 10 10 11 10 16 17 5 7 8 16 22 22 22 22 22 22 22 22 22 22 22 22 22 11 22 16 14 13 15 12 16 
7 1 2 3 20 9 18 9 
5 1 2 20 18 20 
25 1 2 3 9 4 5 6 7 8 9 11 10 16 16 16 22 22 16 22 16 15 13 14 12 16 
4 1 2 18 20 
4 1 2 18 20 
17 1 2 3 20 9 4 6 5 7 8 9 10 10 10 19 17 10 
8 1 2 3 20 9 9 19 9 
24 1 2 20 3 20 9 9 4 5 6 7 8 9 11 10 16 22 22 16 14 12 15 13 16 
4 1 2 18 20 
4 1 2 18 20 
13 1 2 20 3 20 9 9 9 9 9 9 9 19 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 19 9 
5 1 2 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
28 1 2 3 4 6 5 7 8 9 17 5 7 8 10 17 5 7 8 10 17 5 7 8 10 10 17 19 10 
3 1 2 18 
17 1 2 3 20 4 5 6 7 8 9 10 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
15 1 2 3 20 9 4 6 5 7 8 9 10 17 19 10 
8 1 2 3 20 9 9 19 9 
4 1 2 18 20 
5 1 2 20 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
22 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
23 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
31 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 16 16 16 16 13 14 15 12 16 
4 1 2 18 20 
20 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 19 17 10 
24 1 2 3 20 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 18 21 16 
4 1 2 18 20 
5 1 2 20 18 20 
50 1 2 3 20 9 4 5 6 7 8 9 10 10 10 5 17 7 8 10 10 10 10 10 11 10 16 22 22 22 22 22 16 22 22 16 17 5 7 8 16 22 22 22 11 22 14 15 13 12 16 
38 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 11 10 16 16 22 22 22 22 16 22 22 22 13 12 14 15 16 
4 1 2 18 20 
8 1 2 23 23 20 23 18 20 
6 1 2 3 20 18 9 
3 1 2 18 
24 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 16 16 16 16 15 13 12 14 16 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 11 10 18 21 16 
16 1 2 3 9 4 6 5 7 8 9 10 10 10 17 19 10 
20 1 2 3 9 9 4 5 6 7 8 9 10 5 17 7 8 10 19 17 10 
9 1 2 20 3 20 9 9 18 9 
4 1 2 18 20 
25 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 19 17 10 
20 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 16 22 17 19 22 
4 1 2 18 20 
34 1 2 3 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 5 17 7 8 10 11 10 16 18 21 16 
3 1 2 18 
3 1 2 18 
37 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 16 22 16 22 22 22 22 22 22 22 22 13 12 14 15 16 
4 1 2 18 20 
3 1 2 18 
21 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 19 17 22 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 10 11 10 16 16 22 22 14 13 15 12 16 
5 1 2 3 18 9 
24 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 18 21 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 18 21 16 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 11 10 13 15 14 12 16 
8 1 2 20 3 20 9 18 9 
23 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 21 18 16 
5 1 2 3 18 9 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 21 18 16 
23 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 22 22 16 14 12 13 15 16 
23 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 13 14 15 12 16 
3 1 2 18 
8 1 2 3 9 9 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
20 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 19 10 
28 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 17 5 7 8 10 10 10 10 10 19 17 10 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 17 19 10 
3 1 2 18 
24 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 16 14 12 15 13 16 
5 1 2 3 19 9 
6 1 2 3 20 18 9 
5 1 2 3 19 9 
6 1 2 3 20 18 9 
3 1 2 18 
34 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 5 17 7 8 22 22 22 22 22 11 22 16 22 22 14 15 13 12 16 
34 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 11 10 18 21 16 
31 1 2 3 20 9 9 4 5 6 7 8 9 11 10 16 16 22 5 17 7 8 22 22 22 22 22 14 15 13 12 22 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 12 13 15 16 
6 1 2 3 9 19 9 
14 1 2 3 4 5 6 7 8 9 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 17 19 10 
4 1 2 18 20 
22 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 4 9 19 9 
40 1 2 3 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 11 10 5 17 7 8 16 22 22 22 22 22 22 22 11 22 16 15 13 14 12 16 
35 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 16 15 12 13 14 16 
7 1 2 3 20 9 18 9 
33 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 5 17 7 8 16 11 22 13 15 12 14 16 
3 1 2 18 
7 1 2 20 20 20 18 20 
3 1 2 18 
44 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
4 1 2 18 20 
22 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 22 12 15 13 14 16 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
12 1 2 3 4 6 5 7 8 9 17 19 10 
29 1 2 20 3 20 9 4 5 6 7 8 9 11 10 16 22 22 22 22 16 16 22 22 22 15 12 14 13 16 
48 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 11 10 16 16 23 16 16 22 22 22 22 22 22 22 22 16 5 17 7 8 16 14 13 15 12 22 
7 1 2 3 9 4 19 9 
5 1 2 20 18 20 
17 1 2 3 20 9 4 6 5 7 8 9 10 11 10 18 21 16 
17 1 2 3 20 4 6 5 7 8 9 10 11 10 16 21 18 22 
39 1 2 20 20 3 20 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 10 10 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 14 13 12 15 16 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
9 1 2 20 3 20 9 9 19 9 
4 1 2 18 20 
26 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 16 16 14 13 12 15 22 
26 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 16 16 22 22 16 16 14 15 13 12 16 
6 1 2 3 20 18 9 
29 1 2 3 4 5 6 7 8 9 17 5 7 8 10 11 10 16 22 22 5 17 7 8 16 14 15 13 12 22 
33 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 16 22 22 22 14 15 13 12 16 
6 1 2 3 4 18 9 
4 1 2 18 20 
12 1 2 3 4 5 6 7 8 9 19 17 10 
5 1 2 20 18 20 
15 1 2 3 20 9 9 9 9 9 9 9 4 9 19 9 
22 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 18 21 16 
32 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 11 10 16 16 22 16 22 22 22 22 22 22 14 12 13 15 16 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 12 13 15 16 
6 1 2 3 20 18 9 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 10 19 17 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
12 1 2 3 9 9 9 9 9 9 9 19 9 
8 1 2 3 20 9 9 18 9 
18 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 17 19 10 
17 1 2 3 4 6 5 7 8 9 10 10 10 11 10 18 21 16 
5 1 2 3 19 9 
7 1 2 3 20 9 18 9 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
37 1 2 3 20 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 16 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
53 1 2 3 4 5 6 7 8 9 5 17 7 8 10 17 5 7 8 10 10 17 5 7 8 10 10 17 5 7 8 10 10 10 11 10 16 16 22 22 22 22 22 16 5 17 7 8 16 14 12 15 13 22 
17 1 2 3 20 4 5 6 7 8 9 11 10 14 13 12 15 16 
23 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
19 1 2 3 4 6 5 7 8 9 10 11 10 16 22 14 12 13 15 16 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
22 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 
3 1 2 18 
39 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 17 5 7 8 10 17 5 7 8 10 10 10 10 10 10 5 17 7 8 10 17 19 10 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 10 19 17 
9 1 2 3 20 9 9 4 19 9 
26 1 2 3 20 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 
3 1 2 18 
4 1 2 18 20 
26 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 18 21 16 
20 1 2 3 20 9 9 4 5 6 7 8 9 11 10 16 13 15 12 14 16 
36 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 22 22 17 5 7 8 22 22 11 22 14 13 12 15 16 
25 1 2 3 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 18 21 22 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
22 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 19 17 
13 1 2 3 20 4 6 5 7 8 9 17 19 10 
26 1 2 3 20 9 9 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 14 15 13 12 16 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
8 1 2 3 9 9 9 18 9 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 14 13 15 12 16 
14 1 2 3 20 9 4 5 6 7 8 9 17 19 10 
19 1 2 3 4 6 5 7 8 9 10 11 10 16 22 15 14 13 12 16 
3 1 2 18 
21 1 2 3 20 9 9 9 4 5 6 7 8 9 10 11 10 14 13 12 15 16 
10 1 2 3 9 9 9 9 9 9 19 
21 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 12 14 13 15 16 
24 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
17 1 2 3 9 4 6 5 7 8 9 11 10 15 13 14 12 16 
25 1 2 3 20 9 9 4 5 6 7 8 9 11 10 16 16 16 22 22 22 12 15 13 14 16 
3 1 2 18 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
19 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 17 19 10 
6 1 2 3 9 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
28 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 10 19 
5 1 2 3 18 9 
25 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
37 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 11 10 16 14 12 15 13 16 
4 1 2 18 20 
13 1 2 3 9 4 6 5 7 8 9 10 17 19 
3 1 2 18 
13 1 2 3 9 4 5 6 7 8 9 17 19 10 
16 1 2 3 20 9 4 5 6 7 8 9 11 10 21 18 16 
3 1 2 18 
4 1 2 18 20 
34 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 22 22 16 22 22 22 22 22 22 14 13 12 15 16 
38 1 2 20 20 3 20 9 9 9 9 9 9 9 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 16 22 22 22 22 14 12 13 15 16 
14 1 2 3 4 6 5 7 8 9 10 10 19 17 10 
19 1 2 3 20 4 6 5 7 8 9 10 17 5 7 8 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
31 1 2 20 20 20 20 3 20 4 5 6 7 8 9 10 11 10 16 22 22 16 22 16 16 16 22 13 14 12 15 16 
65 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 4 9 9 9 5 6 7 8 9 10 10 10 11 10 16 16 16 16 16 16 22 22 22 22 22 22 22 16 22 22 22 22 16 22 22 22 22 22 22 16 16 16 16 16 16 14 13 12 15 16 
11 1 2 20 3 20 9 9 9 9 9 19 
4 1 2 18 20 
12 1 2 20 3 20 9 9 9 9 9 18 9 
3 1 2 18 
11 1 2 3 9 9 9 9 9 9 9 19 
26 1 2 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 14 15 13 12 16 
28 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 11 10 16 22 22 22 19 17 22 
6 1 2 3 4 19 9 
31 1 2 3 4 5 6 7 8 9 11 10 16 16 16 22 5 17 7 8 22 22 22 22 22 11 22 14 13 12 15 16 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 15 13 12 14 16 
31 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 21 18 16 
11 1 2 3 9 9 9 9 9 9 18 9 
11 1 2 20 3 20 9 9 9 9 18 9 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
29 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 16 22 22 22 22 22 22 19 17 22 
19 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 17 19 10 
6 1 2 3 9 19 9 
5 1 2 20 18 20 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
30 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 11 10 17 5 7 8 16 22 11 22 13 12 14 15 16 
39 1 2 3 20 9 9 9 4 9 5 6 7 8 9 5 17 7 8 10 10 5 17 7 8 10 10 10 11 10 16 16 22 22 22 22 22 18 21 16 
28 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 11 10 16 22 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
30 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 13 14 15 12 22 
21 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
26 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 16 16 22 22 22 22 22 18 21 16 
11 1 2 3 9 9 9 9 9 9 18 9 
25 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 14 13 15 12 22 
4 1 2 18 20 
34 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 17 5 7 8 10 10 11 10 16 22 22 22 14 13 12 15 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
28 1 2 3 4 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 17 5 7 8 10 10 17 19 10 
32 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 11 10 16 22 22 22 22 17 5 7 8 16 15 13 12 14 22 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
5 1 2 23 18 23 
23 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 21 18 22 
5 1 2 3 18 9 
25 1 2 3 9 9 4 6 5 7 8 9 10 10 5 17 7 8 10 11 10 14 13 12 15 16 
34 1 2 3 20 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 21 18 22 
14 1 2 3 9 9 4 5 6 7 8 9 17 19 10 
3 1 2 18 
30 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 17 5 7 8 10 10 10 10 11 10 15 12 13 14 16 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 21 18 16 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
62 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 17 5 7 8 22 17 5 7 8 22 22 22 11 22 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 14 13 15 12 16 
24 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 15 14 12 13 16 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
5 1 2 20 18 20 
21 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 19 
23 1 2 3 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 18 21 16 
27 1 2 20 3 20 9 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 14 15 13 12 16 
3 1 2 18 
30 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 17 5 7 8 16 11 22 13 12 14 15 16 
20 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 14 13 12 15 16 
48 1 2 3 9 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 17 5 7 8 22 22 22 22 22 22 11 22 16 16 16 16 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 19 17 10 
29 1 2 3 20 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 10 17 19 
42 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 17 5 7 8 10 10 11 10 16 22 22 22 22 22 22 22 22 21 18 16 
8 1 2 3 9 9 4 18 9 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 16 16 21 18 16 
8 1 2 3 20 9 9 19 9 
17 1 2 3 9 4 6 5 7 8 9 10 10 11 10 21 18 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 9 9 9 9 4 5 6 7 8 9 11 10 15 14 12 13 16 
3 1 2 18 
19 1 2 3 20 4 5 6 7 8 9 11 10 16 16 14 12 13 15 16 
7 1 2 20 3 20 18 9 
23 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 19 17 10 
33 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 21 18 16 
31 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 19 17 
6 1 2 3 20 18 9 
6 1 2 3 20 18 9 
3 1 2 18 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 9 
51 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 9 9 9 10 9 10 9 9 9 9 9 10 10 10 10 10 10 10 10 10 10 19 17 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 12 13 15 16 
3 1 2 18 
41 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 5 17 7 8 10 10 10 10 11 10 16 22 22 22 5 17 7 8 16 14 13 12 15 22 
22 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 14 12 13 15 16 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 19 17 10 
5 1 2 20 18 20 
3 1 2 18 
5 1 2 20 18 20 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
43 1 2 3 4 5 6 7 8 9 17 5 7 8 10 5 17 7 8 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 19 17 22 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 13 14 12 15 16 
28 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 10 
21 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 11 10 21 18 16 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
25 1 2 3 20 9 9 4 9 5 6 7 8 9 10 10 11 10 16 22 22 14 15 13 12 16 
3 1 2 18 
20 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 16 21 18 16 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
20 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 15 12 14 13 16 
4 1 2 18 20 
22 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 22 18 21 22 
3 1 2 18 
26 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 
4 1 2 18 20 
3 1 2 18 
5 1 2 3 19 9 
22 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 17 5 7 8 10 10 10 
7 1 2 3 20 9 18 9 
5 1 2 3 19 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
5 1 2 20 18 20 
4 1 2 18 20 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 15 13 14 12 16 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
9 1 2 3 9 4 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
29 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 16 16 22 22 22 15 13 12 14 16 
18 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 19 10 17 
19 1 2 3 9 9 4 5 6 7 8 9 10 11 10 14 15 13 12 16 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 17 19 22 
3 1 2 18 
5 1 2 3 19 9 
3 1 2 18 
48 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 23 23 16 16 22 22 5 17 7 8 22 22 22 22 22 22 22 22 22 22 22 11 22 12 13 15 14 16 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
19 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 22 18 21 22 
4 1 2 18 20 
6 1 2 3 20 18 9 
30 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 21 18 16 
3 1 2 18 
27 1 2 3 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 21 18 16 
28 1 2 20 3 20 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 15 12 14 13 16 
18 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
20 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 13 14 12 15 16 
21 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
6 1 2 20 20 18 20 
31 1 2 3 9 4 5 6 7 8 9 11 10 16 22 17 5 7 8 22 22 22 11 22 16 22 22 14 13 15 12 16 
13 1 2 3 20 9 9 9 9 9 9 9 9 19 
3 1 2 18 
45 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 5 17 7 8 10 10 5 17 7 8 10 10 11 10 16 22 22 22 22 22 22 22 19 17 22 
38 1 2 20 3 20 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 11 10 17 5 7 8 16 22 22 22 11 22 16 13 14 12 15 16 
17 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 19 
40 1 2 3 9 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 16 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 19 17 22 
3 1 2 18 
26 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 19 17 10 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 21 18 16 
6 1 2 3 20 19 9 
29 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 16 22 22 22 16 14 12 15 13 16 
20 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
25 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 5 17 7 8 10 10 11 10 
30 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 16 18 21 16 
27 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
6 1 2 3 20 19 9 
45 1 2 3 20 9 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 16 16 22 22 22 16 16 16 22 22 22 22 22 
4 1 2 18 20 
25 1 2 3 20 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 16 13 14 15 12 16 
26 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
7 1 2 3 20 9 18 9 
3 1 2 18 
23 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 11 10 16 12 13 15 14 16 
9 1 2 3 9 9 9 9 19 9 
16 1 2 3 9 4 6 5 7 8 9 10 10 10 10 17 19 
16 1 2 3 4 5 6 7 8 9 10 10 11 10 21 18 16 
34 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 5 17 7 8 10 11 10 16 16 22 22 22 16 16 16 18 21 16 
3 1 2 18 
3 1 2 18 
21 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 19 17 
23 1 2 3 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 19 17 10 
4 1 2 18 20 
32 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 21 18 16 
27 1 2 3 4 9 6 5 7 8 9 5 17 7 8 10 5 17 7 8 10 10 10 10 10 17 19 10 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 11 10 21 18 16 
20 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 15 13 12 14 16 
34 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 16 16 17 5 7 8 16 11 22 14 13 12 15 16 
34 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 16 16 22 22 22 22 22 22 22 22 22 22 16 22 22 22 
17 1 2 3 9 4 6 5 7 8 9 11 10 15 13 12 14 16 
23 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 14 12 13 15 16 
3 1 2 18 
9 1 2 3 20 9 9 9 18 9 
21 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 14 13 15 12 16 
5 1 2 3 19 9 
31 1 2 3 20 4 6 5 7 8 9 11 10 16 16 16 22 22 22 22 22 16 22 22 22 22 22 14 12 13 15 16 
9 1 2 3 9 9 9 9 9 19 
24 1 2 3 4 9 5 6 7 8 9 10 11 10 16 22 22 22 22 22 15 13 12 14 16 
15 1 2 20 3 20 4 6 5 7 8 9 10 19 17 10 
13 1 2 3 4 6 5 7 8 9 10 17 19 10 
29 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
26 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
8 1 2 3 20 9 9 19 9 
26 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 22 22 16 22 22 22 15 13 14 12 16 
4 1 2 18 20 
14 1 2 20 3 20 4 5 6 7 8 9 19 17 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 18 9 
3 1 2 18 
26 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 19 17 
24 1 2 20 20 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 17 19 10 
19 1 2 3 4 5 6 7 8 9 10 10 11 10 16 14 15 13 12 16 
23 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 11 10 16 16 21 18 16 
5 1 2 3 18 9 
21 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 18 21 16 
45 1 2 3 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 5 17 7 8 10 10 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 16 13 14 12 15 16 
4 1 2 18 20 
44 1 2 3 4 5 6 7 8 9 17 5 7 8 10 5 17 7 8 10 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 22 17 5 7 8 22 22 17 19 22 
25 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 12 13 14 15 16 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 19 17 10 
13 1 2 3 9 4 6 5 7 8 9 19 17 10 
29 1 2 3 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 19 17 
7 1 2 3 20 9 18 9 
3 1 2 18 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
20 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
8 1 2 20 3 20 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 19 17 10 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 
23 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 14 15 12 13 16 
26 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
21 1 2 20 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
23 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
33 1 2 3 9 4 5 6 7 8 9 11 10 16 5 17 7 8 16 22 22 22 22 22 22 22 22 11 22 14 12 15 13 16 
12 1 2 3 4 6 5 7 8 9 17 19 10 
6 1 2 20 20 18 20 
4 1 2 18 20 
19 1 2 3 20 9 9 4 6 5 7 8 9 10 11 10 16 19 17 22 
4 1 2 18 20 
19 1 2 3 20 4 6 5 7 8 9 11 10 16 22 15 14 12 13 16 
26 1 2 3 20 4 6 5 7 8 9 10 10 10 5 17 7 8 10 10 10 10 11 10 21 18 16 
24 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 22 14 15 13 12 16 
20 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 22 22 21 18 22 
7 1 2 3 20 9 19 9 
32 1 2 3 4 6 5 7 8 9 11 10 16 16 22 22 16 16 22 22 22 16 22 22 22 22 22 16 14 15 13 12 16 
43 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 22 22 22 16 16 22 22 22 22 22 22 22 22 22 22 16 16 16 16 16 16 16 16 14 12 13 15 16 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 20 9 18 9 
12 1 2 3 9 9 9 9 9 9 9 9 19 
21 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 22 14 15 13 12 16 
7 1 2 3 20 9 18 9 
15 1 2 3 4 6 5 7 8 9 10 10 10 19 17 10 
23 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 16 22 22 12 14 13 15 16 
16 1 2 3 4 6 5 7 8 9 11 10 14 13 15 12 16 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 14 12 15 13 16 
14 1 2 3 9 9 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
17 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 17 19 
5 1 2 3 19 9 
47 1 2 3 20 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 17 5 7 8 16 12 13 14 15 22 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 14 13 12 15 16 
3 1 2 18 
30 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 5 17 7 8 16 14 12 13 15 22 
5 1 2 3 19 9 
3 1 2 18 
26 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 16 16 22 22 22 22 22 19 17 22 
12 1 2 3 20 9 9 9 9 9 9 19 9 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
26 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 16 16 22 22 22 22 13 14 15 12 16 
22 1 2 3 9 9 9 4 6 5 7 8 9 10 10 11 10 16 14 12 13 15 16 
14 1 2 3 4 5 6 7 8 9 11 10 21 18 16 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 19 9 
28 1 2 3 20 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 10 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
41 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 5 17 7 8 10 10 10 10 11 10 16 16 22 22 22 22 16 12 13 15 14 16 
29 1 2 3 20 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
4 1 2 18 20 
29 1 2 3 4 6 5 7 8 9 17 5 7 8 10 5 17 7 8 10 10 5 17 7 8 10 10 17 19 10 
26 1 2 3 9 9 4 5 6 7 8 9 10 10 10 17 5 7 8 10 10 10 10 10 10 17 19 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
19 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 13 15 14 12 16 
19 1 2 3 9 9 9 4 6 5 7 8 9 10 10 11 10 21 18 16 
17 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 
3 1 2 18 
26 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 15 12 14 13 16 
3 1 2 18 
48 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 5 17 7 8 16 22 22 22 22 11 22 13 12 14 15 16 
3 1 2 18 
15 1 2 3 4 6 5 7 8 9 10 11 10 21 18 16 
24 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 14 13 12 15 16 
21 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 13 15 12 14 16 
3 1 2 18 
25 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 16 16 22 22 22 14 13 12 15 16 
23 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 17 5 7 8 10 10 10 
6 1 2 3 20 18 9 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 17 19 
45 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 16 22 22 22 16 16 16 22 22 22 22 17 5 7 8 16 22 22 22 22 11 22 16 16 14 13 12 15 16 
5 1 2 3 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
24 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
17 1 2 3 9 9 9 9 9 4 5 6 7 8 9 17 19 10 
15 1 2 20 3 20 4 6 5 7 8 9 10 19 17 10 
3 1 2 18 
5 1 2 20 18 20 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
5 1 2 3 19 9 
4 1 2 18 20 
4 1 2 18 20 
15 1 2 3 4 6 5 7 8 9 10 10 10 10 19 17 
3 1 2 18 
21 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 10 17 19 10 
12 1 2 3 4 5 6 7 8 9 19 17 10 
6 1 2 3 4 18 9 
4 1 2 18 20 
32 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 22 16 16 16 22 22 13 14 12 15 16 
28 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 17 5 7 8 10 10 10 10 10 10 
4 1 2 18 20 
17 1 2 3 9 4 5 6 7 8 9 10 10 11 10 18 21 16 
4 1 2 18 20 
25 1 2 3 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 14 13 12 15 16 
21 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 17 19 10 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
11 1 2 3 9 9 9 4 9 9 19 9 
16 1 2 3 20 9 9 4 6 5 7 8 9 10 19 17 10 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 18 21 16 
6 1 2 3 9 18 9 
3 1 2 18 
11 1 2 3 20 9 9 9 9 9 18 9 
5 1 2 3 19 9 
22 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 21 18 16 
4 1 2 18 20 
6 1 2 23 23 18 23 
14 1 2 20 3 20 9 4 9 9 9 9 9 19 9 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 18 21 16 
21 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 22 15 13 12 14 16 
7 1 2 3 9 9 19 9 
5 1 2 3 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
23 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 14 12 15 13 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 20 18 9 
43 1 2 3 20 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 16 16 22 22 22 16 22 22 22 22 22 16 16 22 19 17 22 
10 1 2 3 9 9 9 9 9 19 9 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
8 1 2 3 20 9 9 9 19 
26 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
3 1 2 18 
15 1 2 3 9 4 5 6 7 8 9 10 10 10 19 17 
26 1 2 3 4 6 5 7 8 9 11 10 16 22 22 16 22 22 22 22 16 16 14 15 12 13 16 
4 1 2 18 20 
4 1 2 18 20 
6 1 2 3 9 18 9 
6 1 2 3 20 18 9 
17 1 2 3 9 4 5 6 7 8 9 10 10 11 10 18 21 16 
24 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 14 13 15 12 16 
32 1 2 3 20 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 10 10 10 10 5 17 7 8 10 10 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
30 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 10 10 5 17 7 8 10 11 10 14 12 13 15 16 
29 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 16 22 22 22 13 14 15 12 16 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 13 12 15 16 
19 1 2 3 4 6 5 7 8 9 10 10 10 11 10 12 13 14 15 16 
32 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 16 16 16 16 16 16 16 16 12 14 13 15 16 
24 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 17 19 
9 1 2 3 9 9 9 9 9 19 
3 1 2 18 
8 1 2 3 9 9 9 19 9 
21 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 16 22 22 21 18 16 
26 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 14 12 13 15 16 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 18 21 16 
40 1 2 3 20 9 4 5 6 7 8 9 5 17 7 8 10 11 10 16 22 22 16 22 22 22 22 22 22 17 5 7 8 16 11 22 12 14 13 15 16 
3 1 2 18 
7 1 2 3 9 4 18 9 
4 1 2 18 20 
3 1 2 18 
33 1 2 20 3 20 9 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 11 10 21 18 16 
4 1 2 18 20 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 15 13 12 16 
3 1 2 18 
6 1 2 3 9 19 9 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 19 9 
11 1 2 3 20 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
17 1 2 3 20 4 5 6 7 8 9 11 10 14 15 13 12 16 
5 1 2 3 18 9 
26 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 11 10 16 15 13 14 12 16 
3 1 2 18 
27 1 2 3 20 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 5 17 7 8 10 10 11 10 
17 1 2 3 4 5 6 7 8 9 10 11 10 13 12 15 14 16 
18 1 2 20 20 3 20 4 5 6 7 8 9 10 11 10 18 21 16 
27 1 2 20 20 3 20 4 5 6 7 8 9 10 10 10 11 10 16 16 16 16 16 15 13 12 14 16 
18 1 2 3 4 6 5 7 8 9 10 10 11 10 14 12 13 15 16 
27 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 22 14 13 12 15 16 
19 1 2 3 4 6 5 7 8 9 11 10 16 22 16 12 14 13 15 16 
53 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 16 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 
8 1 2 3 9 9 9 9 19 
16 1 2 20 3 20 9 9 9 9 9 9 9 9 9 18 9 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 19 17 
20 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 17 19 
28 1 2 3 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 14 13 15 12 16 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 14 12 13 15 16 
23 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 11 10 14 13 12 15 16 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 10 10 19 17 10 
3 1 2 18 
15 1 2 3 9 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 19 9 
19 1 2 3 20 9 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 12 14 13 15 16 
3 1 2 18 
4 1 2 18 20 
44 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 21 18 16 
12 1 2 3 4 5 6 7 8 9 19 17 10 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 21 18 16 
22 1 2 20 3 20 9 9 9 4 5 6 7 8 9 10 11 10 13 14 15 12 16 
4 1 2 18 20 
9 1 2 3 20 9 9 4 18 9 
24 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 11 10 18 21 16 
23 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 14 13 15 12 16 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
12 1 2 20 3 20 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 20 18 20 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 20 9 19 9 
3 1 2 18 
3 1 2 18 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 19 9 
6 1 2 3 9 18 9 
22 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 11 10 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
10 1 2 20 3 20 9 9 9 18 9 
47 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 22 17 19 22 
29 1 2 3 4 5 6 7 8 9 10 11 10 16 5 17 7 8 22 22 22 22 22 11 22 13 14 12 15 16 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 4 19 9 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 21 18 16 
31 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 15 13 12 16 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
25 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 21 18 10 
3 1 2 18 
40 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 16 16 16 16 16 22 22 16 22 22 22 22 22 16 22 22 22 22 22 16 13 14 15 12 16 
6 1 2 23 23 18 23 
46 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 10 17 5 7 8 10 10 10 11 10 16 22 22 22 22 22 5 17 7 8 22 5 17 7 8 22 22 19 17 22 
3 1 2 18 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 16 13 14 12 15 16 
16 1 2 3 4 6 5 7 8 9 11 10 13 14 12 15 16 
38 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 16 17 5 7 8 22 22 22 17 5 7 8 22 22 22 11 22 13 14 15 12 16 
26 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 15 12 14 13 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 18 9 
23 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 16 22 16 14 12 15 13 16 
5 1 2 3 19 9 
3 1 2 18 
3 1 2 18 
19 1 2 3 9 9 4 6 5 7 8 9 10 11 10 12 15 13 14 16 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
7 1 2 3 9 9 19 9 
25 1 2 20 20 20 20 20 3 20 9 9 4 6 5 7 8 9 10 10 10 11 10 18 21 16 
6 1 2 3 20 18 9 
21 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
6 1 2 3 20 18 9 
3 1 2 18 
5 1 2 20 18 20 
22 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 14 13 12 15 22 
27 1 2 3 9 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 11 10 16 17 19 22 
3 1 2 18 
11 1 2 3 9 9 9 9 9 9 9 19 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 11 10 
19 1 2 3 9 4 6 5 7 8 9 10 10 11 10 14 13 15 12 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
23 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 16 21 18 22 
4 1 2 18 20 
33 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 22 16 17 5 7 8 16 22 22 22 11 22 13 14 15 12 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
5 1 2 3 18 9 
29 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 10 
3 1 2 18 
27 1 2 3 9 9 9 4 6 5 7 8 9 10 10 5 17 7 8 10 10 11 10 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
27 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 14 12 13 15 16 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
7 1 2 20 3 20 18 9 
29 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 5 17 7 8 16 14 15 13 12 22 
21 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 19 17 10 
15 1 2 3 4 6 5 7 8 9 10 10 10 10 17 19 
22 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 18 21 16 
26 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
6 1 2 3 9 19 9 
3 1 2 18 
27 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 15 13 14 12 16 
19 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 19 17 10 
12 1 2 3 4 5 6 7 8 9 19 17 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
14 1 2 3 9 4 5 6 7 8 9 10 19 17 10 
36 1 2 3 9 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 11 10 16 16 22 22 22 22 16 22 16 16 14 13 12 15 16 
4 1 2 18 20 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 16 14 12 15 13 16 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
22 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
20 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 21 18 16 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 17 19 10 
6 1 2 3 9 18 9 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 17 19 10 
4 1 2 18 20 
5 1 2 20 18 20 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 19 9 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 16 22 22 22 21 18 16 
11 1 2 3 9 9 9 9 9 9 9 19 
16 1 2 3 4 5 6 7 8 9 11 10 13 14 15 12 16 
3 1 2 18 
47 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 5 17 7 8 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 16 22 22 17 5 7 8 16 14 13 12 15 22 
3 1 2 18 
27 1 2 3 9 9 9 9 9 4 6 5 7 8 9 11 10 16 22 22 22 16 16 13 15 12 14 16 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 13 14 15 12 16 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 20 20 20 3 20 4 6 5 7 8 9 10 10 10 10 10 19 17 
3 1 2 18 
3 1 2 18 
14 1 2 3 9 9 4 5 6 7 8 9 17 19 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
23 1 2 3 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 11 10 18 21 16 
6 1 2 3 9 18 9 
3 1 2 18 
3 1 2 18 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 17 19 
4 1 2 18 20 
7 1 2 20 20 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
14 1 2 3 9 4 6 5 7 8 9 10 18 21 10 
23 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
30 1 2 20 3 20 4 5 6 7 8 9 10 17 5 7 8 10 17 5 7 8 10 10 10 10 10 10 19 17 10 
16 1 2 3 20 4 6 5 7 8 9 10 11 10 18 21 16 
5 1 2 20 18 20 
16 1 2 3 20 9 4 5 6 7 8 9 11 10 21 18 16 
3 1 2 18 
3 1 2 18 
22 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 19 17 
7 1 2 3 9 9 18 9 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
17 1 2 3 4 6 5 7 8 9 10 10 10 10 10 17 19 10 
3 1 2 18 
22 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 19 
10 1 2 3 9 9 9 9 9 19 9 
7 1 2 3 20 9 18 9 
3 1 2 18 
14 1 2 3 20 4 5 6 7 8 9 10 19 17 10 
9 1 2 3 9 9 9 9 18 9 
32 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 22 22 22 16 22 22 22 22 22 22 21 18 16 
4 1 2 18 20 
9 1 2 3 9 9 9 9 18 9 
16 1 2 3 9 4 6 5 7 8 9 10 10 10 10 19 17 
3 1 2 18 
12 1 2 3 9 9 9 9 9 9 9 19 9 
25 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 
29 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 16 14 13 15 12 16 
23 1 2 3 4 6 5 7 8 9 11 10 16 22 22 16 22 22 16 13 14 15 12 16 
8 1 2 3 9 9 9 18 9 
4 1 2 18 20 
27 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 10 19 17 
30 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 5 17 7 8 22 22 22 22 17 19 22 
14 1 2 20 3 20 4 5 6 7 8 9 19 17 10 
4 1 2 18 20 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
34 1 2 3 9 9 4 9 6 5 7 8 9 10 17 5 7 8 10 10 10 10 10 11 10 16 16 16 22 22 22 22 21 18 22 
6 1 2 20 20 18 20 
5 1 2 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
22 1 2 20 3 20 9 9 4 6 5 7 8 9 10 10 11 10 14 13 12 15 16 
3 1 2 18 
26 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 17 19 10 
12 1 2 3 9 9 9 9 9 9 9 19 9 
7 1 2 20 3 20 18 9 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
42 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 16 16 22 22 22 22 22 22 22 22 22 22 22 22 16 22 22 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
22 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 11 10 13 14 12 15 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 17 19 10 
23 1 2 20 3 20 9 4 5 6 7 8 9 10 17 5 7 8 10 11 10 18 21 16 
24 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 17 5 7 8 10 18 21 10 
21 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 19 17 10 
4 1 2 18 20 
8 1 2 3 9 9 9 19 9 
20 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 21 18 10 
4 1 2 18 20 
25 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
37 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 11 10 16 22 22 22 16 22 22 16 5 17 7 8 16 12 14 15 13 22 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
5 1 2 3 19 9 
26 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 16 22 22 14 12 13 15 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 17 5 7 8 10 10 10 
3 1 2 18 
18 1 2 20 3 20 9 9 9 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
11 1 2 3 20 9 9 9 9 9 18 9 
24 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 19 17 
23 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 19 17 
3 1 2 18 
5 1 2 3 19 9 
7 1 2 3 9 4 19 9 
7 1 2 20 3 20 18 9 
7 1 2 3 20 9 19 9 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
17 1 2 3 9 4 6 5 7 8 9 10 10 11 10 18 21 16 
4 1 2 18 20 
4 1 2 18 20 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
20 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 10 10 17 19 
31 1 2 3 20 9 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 10 10 10 17 19 
23 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 22 16 15 12 13 14 16 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 16 16 16 22 22 17 19 22 
14 1 2 3 4 5 6 7 8 9 11 10 18 21 16 
3 1 2 18 
7 1 2 3 20 9 18 9 
5 1 2 3 18 9 
7 1 2 3 20 9 18 9 
21 1 2 3 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 17 19 10 
44 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 22 11 22 14 13 12 15 16 
27 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 21 18 22 
8 1 2 3 9 9 9 19 9 
4 1 2 18 20 
34 1 2 3 9 9 4 9 9 5 6 7 8 9 5 17 7 8 10 5 17 7 8 10 17 5 7 8 10 10 10 10 17 19 10 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 13 14 15 12 16 
12 1 2 3 4 5 6 7 8 9 19 17 10 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 19 9 
5 1 2 3 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 10 10 18 21 10 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 
24 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 
35 1 2 3 20 9 9 9 4 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 10 10 10 10 11 10 16 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
32 1 2 3 20 9 4 6 5 7 8 9 10 10 11 10 16 16 16 22 22 22 22 22 22 22 16 16 14 12 13 15 16 
6 1 2 3 9 18 9 
47 1 2 3 20 4 5 6 7 8 9 10 10 17 5 7 8 10 11 10 16 16 16 22 22 22 22 17 5 7 8 22 22 22 22 22 11 22 16 16 22 22 22 14 13 12 15 16 
26 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 11 10 16 22 22 14 15 13 12 16 
6 1 2 3 9 18 9 
4 1 2 18 20 
29 1 2 20 20 20 3 20 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 11 10 16 18 21 16 
31 1 2 3 9 9 9 9 9 9 9 9 4 6 5 7 8 9 11 10 16 22 22 22 22 16 16 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
13 1 2 3 4 6 5 7 8 9 10 18 21 10 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 9 9 4 5 6 7 8 9 11 10 16 22 22 16 14 15 12 13 16 
3 1 2 18 
3 1 2 18 
10 1 2 3 20 9 9 9 9 18 9 
32 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 16 16 16 16 16 22 22 14 12 13 15 16 
44 1 2 3 20 4 6 5 7 8 9 5 17 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 16 14 12 13 15 16 
4 1 2 18 20 
3 1 2 18 
26 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 12 14 15 13 16 
40 1 2 3 4 6 5 7 8 9 10 10 10 11 10 5 17 7 8 16 22 22 11 22 16 16 22 22 22 22 22 22 16 16 16 16 14 15 12 13 16 
7 1 2 3 20 9 19 9 
23 1 2 20 20 20 3 20 9 9 4 5 6 7 8 9 10 11 10 13 14 15 12 16 
7 1 2 3 20 9 18 9 
42 1 2 3 20 9 9 4 9 9 9 9 9 9 6 5 7 8 9 11 10 16 22 22 22 22 22 22 16 16 22 5 17 7 8 22 22 22 12 14 13 15 22 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
5 1 2 3 18 9 
3 1 2 18 
10 1 2 3 9 9 9 9 4 19 9 
6 1 2 3 20 18 9 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 18 9 
31 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 22 22 16 22 22 22 22 14 15 12 13 22 
22 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
6 1 2 3 9 19 9 
3 1 2 18 
24 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 16 16 18 21 16 
40 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 10 10 11 10 16 16 22 22 22 22 5 17 7 8 16 14 12 13 15 22 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 13 12 14 15 16 
11 1 2 3 20 9 9 9 9 9 18 9 
21 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 21 18 10 
4 1 2 18 20 
37 1 2 20 3 20 9 9 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 10 10 10 10 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
29 1 2 3 4 5 6 7 8 9 10 10 11 10 5 17 7 8 16 22 22 22 22 11 22 13 12 14 15 16 
18 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 19 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
19 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 19 17 10 
19 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 18 21 10 
4 1 2 18 20 
3 1 2 18 
8 1 2 3 9 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
5 1 2 20 18 20 
32 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 16 22 22 22 22 22 22 22 22 19 17 22 
11 1 2 3 4 9 9 9 9 9 19 9 
8 1 2 3 9 9 9 19 9 
5 1 2 20 18 20 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 9 18 9 
4 1 2 18 20 
3 1 2 18 
36 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 22 16 22 22 22 22 22 22 16 12 15 14 13 16 
5 1 2 3 18 9 
24 1 2 20 3 20 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 18 21 16 
5 1 2 20 18 20 
25 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 14 13 12 15 16 
6 1 2 3 9 19 9 
4 1 2 18 20 
33 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 21 18 22 
6 1 2 3 20 18 9 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 19 17 
17 1 2 3 4 5 6 7 8 9 5 17 7 8 10 19 17 10 
8 1 2 3 9 9 9 19 9 
9 1 2 3 9 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 19 17 10 
3 1 2 18 
20 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
23 1 2 3 4 9 6 5 7 8 9 10 10 10 11 10 16 16 16 15 13 14 12 16 
4 1 2 18 20 
21 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 21 18 16 
32 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 11 10 16 17 5 7 8 16 14 12 15 13 22 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 17 19 10 
24 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
28 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 5 17 7 8 10 11 10 12 14 13 15 16 
3 1 2 18 
30 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 13 12 14 15 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
8 1 2 3 9 9 9 19 9 
4 1 2 18 20 
18 1 2 3 4 6 5 7 8 9 11 10 16 22 13 14 15 12 16 
22 1 2 3 20 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 
4 1 2 18 20 
3 1 2 18 
23 1 2 3 20 9 4 5 6 7 8 9 10 10 10 10 10 5 17 7 8 10 10 10 
3 1 2 18 
9 1 2 3 9 9 9 9 18 9 
15 1 2 3 4 6 5 7 8 9 10 11 10 21 18 16 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
22 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 21 18 16 
19 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
34 1 2 3 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 11 10 16 22 22 22 22 22 22 16 16 22 17 19 22 
10 1 2 3 9 9 9 9 4 19 9 
31 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 16 16 13 14 15 12 16 
7 1 2 3 20 4 18 9 
4 1 2 18 20 
55 1 2 3 20 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 5 17 7 8 22 22 22 22 17 5 7 8 22 22 22 5 17 7 8 22 22 22 22 11 22 16 14 15 12 13 16 
26 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 12 13 15 14 16 
18 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 
23 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
3 1 2 18 
9 1 2 3 20 9 9 9 19 9 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 18 21 16 
14 1 2 3 9 9 4 5 6 7 8 9 10 10 10 
24 1 2 3 20 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 15 13 12 14 16 
3 1 2 18 
3 1 2 18 
38 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 16 16 16 22 22 16 22 22 22 22 14 12 15 13 16 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 9 19 9 
42 1 2 3 4 5 6 7 8 9 17 5 7 8 10 17 5 7 8 10 10 10 10 10 10 11 10 16 16 22 22 22 22 16 22 16 16 16 14 15 12 13 16 
17 1 2 3 9 9 9 9 4 5 6 7 8 9 10 19 17 10 
3 1 2 18 
6 1 2 3 20 19 9 
26 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 
19 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 17 19 10 
5 1 2 3 18 9 
12 1 2 3 4 6 5 7 8 9 19 17 10 
29 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 15 12 14 13 16 
3 1 2 18 
55 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 16 16 22 22 5 17 7 8 22 22 5 17 7 8 22 17 5 7 8 22 22 22 11 22 14 13 12 15 16 
22 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 
29 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 16 22 15 14 12 13 16 
4 1 2 18 20 
49 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 5 7 8 10 10 10 11 10 16 22 22 22 22 16 22 22 16 22 22 22 16 12 14 15 13 16 
9 1 2 3 20 9 9 9 19 9 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 
32 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 16 22 22 22 22 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
21 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 5 17 7 8 10 10 
30 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 17 5 7 8 10 10 11 10 14 12 13 15 16 
17 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 10 
21 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 
3 1 2 18 
24 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 18 21 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
26 1 2 3 20 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 16 13 12 14 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 9 18 9 
5 1 2 20 18 20 
5 1 2 20 18 20 
6 1 2 20 20 18 20 
33 1 2 3 20 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 11 10 16 22 22 22 22 13 14 12 15 16 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
5 1 2 3 19 9 
7 1 2 3 9 9 9 9 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 11 10 14 13 15 12 16 
3 1 2 18 
32 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 11 10 16 16 16 16 16 16 16 22 22 22 22 22 22 22 22 
3 1 2 18 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
8 1 2 3 9 9 9 9 9 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
6 1 2 3 20 18 9 
26 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 22 22 22 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
37 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 13 14 12 15 16 
32 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 5 17 7 8 10 10 10 10 11 10 15 12 13 14 16 
11 1 2 3 9 9 9 9 9 9 9 9 
8 1 2 20 3 20 9 18 9 
3 1 2 18 
17 1 2 20 3 20 4 5 6 7 8 9 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 19 9 
23 1 2 3 20 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 18 21 16 
7 1 2 3 9 9 18 9 
17 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
12 1 2 3 20 9 9 9 9 9 9 18 9 
34 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 22 22 22 22 22 16 16 14 12 15 13 16 
7 1 2 3 9 9 9 9 
7 1 2 3 20 9 19 9 
3 1 2 18 
26 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
24 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 17 5 7 8 10 10 
21 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 
14 1 2 3 9 9 9 4 6 5 7 8 9 10 10 
6 1 2 3 4 19 9 
24 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 11 10 16 22 22 22 
17 1 2 3 4 6 5 7 8 9 11 10 16 22 22 18 21 16 
10 1 2 3 9 9 9 9 9 19 9 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
5 1 2 20 18 20 
5 1 2 23 18 23 
38 1 2 20 20 20 20 20 20 20 3 20 4 5 6 7 8 9 10 10 10 11 10 17 5 7 8 16 22 22 22 22 11 22 15 12 13 14 16 
20 1 2 3 4 6 5 7 8 9 10 10 10 10 11 10 13 15 14 12 16 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
23 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 16 18 21 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 18 21 16 
22 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
7 1 2 20 20 20 18 20 
25 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 14 13 12 15 16 
28 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 16 22 22 18 21 22 
6 1 2 3 20 19 9 
22 1 2 3 20 4 5 6 7 8 9 10 11 10 16 22 22 22 15 14 12 13 16 
4 1 2 18 20 
5 1 2 3 18 9 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
12 1 2 3 20 9 9 9 9 9 9 18 9 
4 1 2 18 20 
10 1 2 20 3 20 9 9 9 19 9 
3 1 2 18 
33 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 16 22 22 22 22 14 13 15 12 16 
35 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 16 17 5 7 8 16 22 22 11 22 14 15 13 12 16 
3 1 2 18 
20 1 2 20 3 20 4 5 6 7 8 9 10 10 10 11 10 16 18 21 16 
15 1 2 20 3 20 4 5 6 7 8 9 10 19 17 10 
29 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 16 22 22 22 22 22 17 19 22 
4 1 2 18 20 
3 1 2 18 
23 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 22 16 16 14 13 15 12 16 
3 1 2 18 
7 1 2 20 20 20 18 20 
31 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 22 22 22 22 22 22 22 16 14 12 13 15 16 
4 1 2 18 20 
3 1 2 18 
7 1 2 20 20 20 18 20 
3 1 2 18 
3 1 2 18 
6 1 2 20 20 18 20 
19 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 
3 1 2 18 
14 1 2 3 9 9 4 5 6 7 8 9 17 19 10 
35 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 16 22 22 22 16 22 22 22 22 22 16 22 22 16 16 22 
22 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 22 14 13 12 15 16 
17 1 2 3 9 4 5 6 7 8 9 10 10 17 5 7 8 10 
8 1 2 3 20 9 9 18 9 
5 1 2 20 18 20 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
23 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
27 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 22 22 13 12 14 15 16 
16 1 2 20 3 20 4 6 5 7 8 9 10 10 17 19 10 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 10 10 10 17 19 10 
4 1 2 18 20 
3 1 2 18 
20 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 14 13 12 15 16 
3 1 2 18 
27 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 11 10 16 22 22 16 16 13 14 15 12 16 
4 1 2 18 20 
14 1 2 3 9 9 4 6 5 7 8 9 10 10 10 
3 1 2 18 
3 1 2 18 
36 1 2 3 20 9 9 4 5 6 7 8 9 10 10 11 10 16 16 16 16 22 22 22 22 22 16 22 22 22 16 16 14 13 15 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 18 9 
23 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 14 13 15 12 16 
21 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 16 16 22 21 18 22 
5 1 2 23 18 23 
3 1 2 18 
25 1 2 3 20 9 4 6 5 7 8 9 17 5 7 8 10 10 5 17 7 8 10 10 10 10 
5 1 2 20 18 20 
4 1 2 18 20 
8 1 2 20 3 20 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 16 22 18 21 22 
5 1 2 20 18 20 
3 1 2 18 
25 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 22 14 12 13 15 16 
3 1 2 18 
10 1 2 3 9 9 9 9 9 18 9 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 10 10 17 19 10 
7 1 2 3 20 9 18 9 
17 1 2 3 9 4 5 6 7 8 9 11 10 15 13 12 14 16 
7 1 2 3 20 9 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 20 4 6 5 7 8 9 10 11 10 14 13 12 15 16 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 10 5 17 7 8 10 10 10 
6 1 2 3 20 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 4 19 9 
3 1 2 18 
23 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 16 22 22 
20 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 
4 1 2 18 20 
31 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 22 22 16 5 17 7 8 16 14 15 13 12 22 
17 1 2 3 4 5 6 7 8 9 10 11 10 15 13 12 14 16 
3 1 2 18 
6 1 2 3 9 19 9 
16 1 2 3 9 4 6 5 7 8 9 10 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
34 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 17 19 22 
4 1 2 18 20 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 15 13 12 14 16 
17 1 2 3 9 4 6 5 7 8 9 11 10 12 14 13 15 16 
3 1 2 18 
3 1 2 18 
5 1 2 3 19 9 
4 1 2 18 20 
20 1 2 3 20 9 9 9 4 6 5 7 8 9 11 10 14 12 13 15 16 
3 1 2 18 
39 1 2 3 20 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 22 22 22 5 17 7 8 22 22 
20 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 17 5 7 8 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
24 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 14 15 13 12 16 
7 1 2 3 9 9 18 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 17 19 10 
21 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 11 10 16 18 21 16 
6 1 2 3 20 19 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
12 1 2 3 4 6 5 7 8 9 19 17 10 
23 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 15 14 12 13 16 
18 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 
16 1 2 3 4 6 5 7 8 9 10 10 11 10 21 18 16 
3 1 2 18 
5 1 2 3 19 9 
4 1 2 18 20 
4 1 2 18 20 
22 1 2 3 4 5 6 7 8 9 10 10 10 11 10 16 22 22 14 12 15 13 16 
12 1 2 3 4 5 6 7 8 9 17 19 10 
21 1 2 3 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 19 17 10 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 18 21 16 
3 1 2 18 
5 1 2 20 18 20 
4 1 2 18 20 
4 1 2 18 20 
29 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 22 22 22 13 14 15 12 16 
18 1 2 3 9 9 4 5 6 7 8 9 11 10 13 12 14 15 16 
5 1 2 20 18 20 
3 1 2 18 
7 1 2 3 9 9 19 9 
26 1 2 3 20 4 5 6 7 8 9 10 10 10 11 10 16 22 22 22 22 22 14 13 12 15 16 
22 1 2 3 20 9 9 9 9 4 5 6 7 8 9 11 10 16 16 16 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
30 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 22 22 16 22 22 22 22 13 14 12 15 16 
3 1 2 18 
26 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 
4 1 2 18 20 
25 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 21 18 22 
5 1 2 20 18 20 
20 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 
16 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
31 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 
42 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 16 16 16 16 22 5 17 7 8 22 22 22 22 22 22 11 22 14 13 12 15 16 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 14 15 12 13 16 
36 1 2 3 20 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 17 5 7 8 10 5 17 7 8 10 10 10 10 10 10 10 10 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 16 18 21 16 
4 1 2 18 20 
4 1 2 18 20 
14 1 2 3 20 4 6 5 7 8 9 10 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
13 1 2 3 9 9 9 9 9 9 9 9 9 9 
60 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 16 16 16 22 22 22 16 16 16 16 22 22 22 22 5 17 7 8 22 13 12 14 15 22 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
22 1 2 3 9 4 5 6 7 8 9 10 5 17 7 8 10 11 10 16 21 18 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
21 1 2 20 3 20 9 4 5 6 7 8 9 10 11 10 16 12 14 13 15 16 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 14 15 13 12 16 
3 1 2 18 
3 1 2 18 
19 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 
3 1 2 18 
44 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 16 22 22 17 5 7 8 22 22 22 22 11 22 16 12 14 13 15 16 
22 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 17 5 7 8 10 10 10 
4 1 2 18 20 
17 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 
44 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 22 22 16 16 16 16 16 16 16 22 22 22 22 16 22 22 22 22 22 16 14 13 15 12 16 
21 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 21 18 16 
8 1 2 3 20 9 9 18 9 
6 1 2 3 20 18 9 
3 1 2 18 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
3 1 2 18 
25 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 11 10 16 22 22 22 
18 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 10 10 10 
3 1 2 18 
6 1 2 3 9 9 9 
7 1 2 3 20 9 19 9 
14 1 2 3 9 4 6 5 7 8 9 10 10 10 10 
3 1 2 18 
34 1 2 3 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 10 5 17 7 8 10 10 11 10 16 22 14 12 13 15 16 
4 1 2 18 20 
24 1 2 3 20 9 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 21 18 16 
42 1 2 3 20 9 9 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 22 22 22 16 16 5 17 7 8 22 22 22 22 22 22 22 22 22 
6 1 2 3 20 18 9 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 16 22 19 17 22 
25 1 2 3 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 18 21 16 
16 1 2 3 4 5 6 7 8 9 10 10 10 10 17 19 10 
15 1 2 3 4 6 5 7 8 9 10 10 10 10 10 10 
4 1 2 18 20 
3 1 2 18 
19 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 
26 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 10 10 10 17 5 7 8 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
15 1 2 3 4 6 5 7 8 9 11 10 16 19 17 22 
4 1 2 18 20 
3 1 2 18 
29 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 16 16 16 22 22 22 22 16 21 18 16 
3 1 2 18 
31 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 16 22 22 22 22 22 22 22 22 22 14 12 13 15 16 
7 1 2 3 9 9 18 9 
3 1 2 18 
24 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 11 10 16 23 14 13 12 15 16 
8 1 2 3 9 9 9 19 9 
4 1 2 18 20 
3 1 2 18 
32 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 17 5 7 8 10 10 11 10 16 22 22 22 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 15 14 12 13 16 
7 1 2 3 9 9 19 9 
10 1 2 20 3 20 9 9 9 18 9 
30 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 17 5 7 8 10 10 10 11 10 16 15 13 12 14 16 
9 1 2 3 9 9 9 9 19 9 
8 1 2 3 9 9 9 18 9 
19 1 2 3 9 9 4 9 6 5 7 8 9 10 10 11 10 21 18 16 
6 1 2 3 20 18 9 
19 1 2 3 9 4 6 5 7 8 9 10 11 10 16 13 12 15 14 16 
6 1 2 3 20 18 9 
11 1 2 3 20 9 9 9 9 9 19 9 
35 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 11 10 5 17 7 8 16 22 22 22 22 22 22 22 22 22 22 22 22 22 
4 1 2 18 20 
14 1 2 3 9 9 4 5 6 7 8 9 17 19 10 
3 1 2 18 
7 1 2 3 9 9 18 9 
12 1 2 3 4 5 6 7 8 9 17 19 10 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 20 9 9 9 4 5 6 7 8 9 10 10 10 17 19 10 
6 1 2 3 20 18 9 
5 1 2 3 18 9 
25 1 2 3 20 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 16 14 13 12 15 16 
3 1 2 18 
39 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 11 10 16 16 16 16 22 22 22 16 16 16 22 22 22 13 14 12 15 16 
3 1 2 18 
3 1 2 18 
25 1 2 3 9 9 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 14 13 12 15 16 
3 1 2 18 
10 1 2 3 9 9 9 9 9 19 9 
19 1 2 20 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 10 
20 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 14 15 13 12 16 
21 1 2 3 20 9 4 6 5 7 8 9 10 10 11 10 16 14 12 13 15 22 
22 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 21 18 16 
13 1 2 3 9 9 9 9 9 9 9 9 9 9 
7 1 2 3 9 9 19 9 
11 1 2 3 20 9 9 9 9 9 18 9 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
14 1 2 3 9 9 4 6 5 7 8 9 19 17 10 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
9 1 2 3 20 9 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
8 1 2 3 9 9 9 19 9 
3 1 2 18 
15 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 
3 1 2 18 
26 1 2 3 9 9 9 9 9 4 6 5 7 8 9 11 10 16 22 22 22 22 14 13 12 15 16 
19 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 
3 1 2 18 
20 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 11 10 19 17 16 
48 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 22 5 17 7 8 22 22 22 22 22 22 22 11 22 14 12 13 15 16 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 9 
4 1 2 18 20 
13 1 2 3 4 6 5 7 8 9 10 17 19 10 
3 1 2 18 
17 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 10 
6 1 2 20 20 18 20 
6 1 2 3 9 19 9 
8 1 2 3 20 9 9 18 9 
18 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 18 21 16 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
4 1 2 18 20 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
7 1 2 3 20 9 18 9 
3 1 2 18 
4 1 2 18 20 
41 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 22 16 16 22 16 22 22 22 16 16 17 5 7 8 22 22 22 22 11 22 14 12 13 15 16 
4 1 2 18 20 
4 1 2 18 20 
21 1 2 3 9 4 6 5 7 8 9 11 10 16 16 16 16 13 14 15 12 16 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
26 1 2 3 20 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 
4 1 2 18 20 
23 1 2 3 20 4 6 5 7 8 9 10 5 17 7 8 10 10 11 10 16 18 21 16 
4 1 2 18 20 
30 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 10 11 10 16 16 22 22 22 14 12 13 15 16 
3 1 2 18 
6 1 2 3 9 18 9 
18 1 2 3 20 4 6 5 7 8 9 10 10 10 10 10 10 10 10 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
7 1 2 3 9 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 19 9 
17 1 2 3 20 4 6 5 7 8 9 10 10 10 10 19 17 10 
17 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 10 10 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 20 18 20 
46 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 17 5 7 8 10 5 17 7 8 10 10 10 10 11 10 16 21 18 16 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 9 9 
3 1 2 18 
5 1 2 3 18 9 
12 1 2 3 9 9 9 9 9 9 9 9 9 
28 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 16 22 22 18 21 16 
7 1 2 3 20 9 19 9 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 20 4 5 6 7 8 9 11 10 16 12 14 13 15 16 
8 1 2 3 20 9 9 18 9 
5 1 2 3 18 9 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
19 1 2 3 9 4 5 6 7 8 9 10 10 11 10 14 13 12 15 16 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 9 9 19 9 
25 1 2 3 20 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 16 13 14 12 15 16 
24 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 10 
3 1 2 18 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 10 10 10 11 10 21 18 16 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 17 19 10 
22 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 11 10 21 18 16 
17 1 2 3 20 9 9 4 5 6 7 8 9 10 10 19 17 10 
15 1 2 3 9 4 5 6 7 8 9 10 10 17 19 10 
7 1 2 3 9 9 19 9 
9 1 2 3 9 9 9 9 9 9 
4 1 2 18 20 
22 1 2 3 9 9 9 9 4 6 5 7 8 9 10 11 10 16 14 13 15 12 16 
21 1 2 3 9 4 6 5 7 8 9 10 10 10 10 11 10 15 14 12 13 16 
13 1 2 3 9 9 9 9 9 9 9 9 9 9 
40 1 2 3 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 16 16 22 22 22 22 22 22 22 5 17 7 8 16 13 14 12 15 22 
12 1 2 3 9 9 9 9 9 9 9 9 9 
3 1 2 18 
3 1 2 18 
19 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 
6 1 2 3 9 18 9 
15 1 2 3 9 9 9 4 5 6 7 8 9 19 17 10 
3 1 2 18 
4 1 2 18 20 
7 1 2 3 9 9 19 9 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
22 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 11 10 12 13 14 15 16 
35 1 2 3 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 16 22 22 22 17 5 7 8 16 12 13 15 14 22 
14 1 2 3 9 9 9 9 4 5 6 7 8 9 10 
16 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 
5 1 2 3 18 9 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 19 17 10 
16 1 2 3 9 9 4 6 5 7 8 9 10 10 17 19 10 
28 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 11 10 16 16 22 22 22 22 12 13 15 14 22 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
23 1 2 3 4 6 5 7 8 9 17 5 7 8 10 11 10 16 16 13 14 15 12 16 
3 1 2 18 
14 1 2 3 20 9 4 6 5 7 8 9 10 10 10 
9 1 2 3 20 9 4 9 19 9 
11 1 2 20 3 20 9 9 9 9 19 9 
5 1 2 20 18 20 
16 1 2 20 3 20 4 5 6 7 8 9 10 10 10 10 10 
40 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 16 5 17 7 8 16 22 22 22 22 22 22 22 22 11 22 16 22 22 22 22 22 16 16 16 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
4 1 2 18 20 
10 1 2 3 20 9 9 9 9 18 9 
4 1 2 18 20 
5 1 2 3 19 9 
34 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 22 22 16 16 22 22 22 22 22 13 14 12 15 22 
22 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 17 5 7 8 10 10 
4 1 2 18 20 
10 1 2 20 20 20 3 20 9 18 9 
15 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 
19 1 2 3 9 4 5 6 7 8 9 10 10 10 10 11 10 21 18 16 
16 1 2 3 4 6 5 7 8 9 11 10 14 15 13 12 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
21 1 2 3 4 5 6 7 8 9 10 10 10 10 10 11 10 14 13 15 12 16 
3 1 2 18 
7 1 2 3 9 9 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
17 1 2 3 4 5 6 7 8 9 11 10 16 14 15 12 13 16 
4 1 2 18 20 
8 1 2 3 20 9 9 19 9 
3 1 2 18 
15 1 2 3 20 4 5 6 7 8 9 11 10 18 21 16 
31 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 16 16 5 17 7 8 16 14 15 13 12 22 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
3 1 2 18 
30 1 2 3 4 9 5 6 7 8 9 10 10 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 19 17 22 
3 1 2 18 
19 1 2 3 20 9 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
13 1 2 3 9 9 9 9 9 9 9 9 9 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
3 1 2 18 
20 1 2 3 4 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 13 14 12 15 16 
4 1 2 18 20 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 9 
21 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 22 14 13 15 12 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 17 19 10 
28 1 2 20 3 20 4 5 6 7 8 9 10 10 10 10 11 10 16 16 22 22 22 22 14 13 15 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
26 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 16 13 14 12 15 16 
14 1 2 23 23 23 20 23 23 23 23 23 23 18 20 
14 1 2 23 23 20 20 23 23 23 23 23 23 18 20 
17 1 2 3 9 4 5 6 7 8 9 11 10 13 14 12 15 16 
17 1 2 3 9 9 4 5 6 7 8 9 10 11 10 19 17 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
21 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 10 10 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 9 
12 1 2 3 4 5 6 7 8 9 10 10 10 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
16 1 2 3 4 6 5 7 8 9 11 10 13 14 15 12 16 
4 1 2 18 20 
25 1 2 3 4 5 6 7 8 9 11 10 5 17 7 8 16 22 22 22 22 22 22 17 19 22 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
9 1 2 3 20 9 9 9 19 9 
18 1 2 20 3 20 9 4 6 5 7 8 9 10 11 10 18 21 16 
12 1 2 3 4 6 5 7 8 9 10 10 10 
33 1 2 3 4 6 5 7 8 9 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 14 15 13 12 16 
13 1 2 3 20 9 9 9 9 9 9 9 9 9 
40 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 17 5 7 8 16 22 22 22 11 22 16 22 22 22 22 16 16 22 16 16 14 13 12 15 16 
11 1 2 3 9 9 9 9 9 9 19 9 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
11 1 2 3 9 4 6 5 7 8 9 10 
9 1 2 3 9 9 9 9 19 9 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 10 11 10 
9 1 2 3 9 9 9 9 19 9 
17 1 2 3 20 9 4 6 5 7 8 9 10 11 10 18 21 16 
3 1 2 18 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 10 10 10 11 10 
24 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 16 16 16 16 22 17 19 22 
13 1 2 3 9 4 5 6 7 8 9 17 19 10 
6 1 2 3 20 18 9 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 9 9 
16 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 
3 1 2 18 
19 1 2 3 9 9 9 4 5 6 7 8 9 11 10 12 15 13 14 16 
16 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 
3 1 2 18 
15 1 2 3 9 4 6 5 7 8 9 11 10 18 21 16 
39 1 2 3 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 16 22 22 22 22 22 5 17 7 8 22 22 22 22 11 22 13 14 12 15 16 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 9 9 19 9 
17 1 2 3 4 6 5 7 8 9 10 11 10 14 13 15 12 16 
7 1 2 3 20 9 19 9 
27 1 2 20 3 20 9 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 14 15 13 12 16 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
17 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 11 10 
44 1 2 3 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 5 17 7 8 10 10 10 11 10 16 22 22 22 22 22 22 16 22 22 14 12 13 15 16 
6 1 2 3 20 18 9 
15 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 
3 1 2 18 
6 1 2 3 9 19 9 
26 1 2 3 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 10 19 17 10 
16 1 2 3 4 5 6 7 8 9 11 10 12 13 15 14 16 
20 1 2 3 20 9 4 5 6 7 8 9 11 10 16 22 22 22 21 18 16 
3 1 2 18 
4 1 2 18 20 
15 1 2 3 20 4 5 6 7 8 9 10 10 10 10 10 
17 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 
6 1 2 3 9 19 9 
4 1 2 18 20 
4 1 2 18 20 
5 1 2 3 19 9 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 17 19 10 
22 1 2 3 9 9 4 5 6 7 8 9 11 10 16 16 22 22 13 14 12 15 16 
18 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 
6 1 2 3 20 18 9 
9 1 2 3 20 9 9 9 18 9 
26 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 17 5 7 8 10 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
6 1 2 3 9 18 9 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 13 14 12 15 16 
21 1 2 20 20 3 20 4 5 6 7 8 9 10 10 11 10 14 13 15 12 16 
5 1 2 20 18 20 
16 1 2 3 4 5 6 7 8 9 10 11 10 16 21 18 22 
3 1 2 18 
22 1 2 3 9 9 9 4 6 5 7 8 9 11 10 16 22 16 14 13 12 15 16 
9 1 2 3 9 9 9 9 19 9 
20 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 
26 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 22 16 16 16 12 13 15 14 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 14 13 12 15 16 
35 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 11 10 16 16 16 5 17 7 8 16 14 13 12 15 22 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 12 13 15 14 16 
14 1 2 3 9 4 6 5 7 8 9 10 10 10 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
25 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 5 17 7 8 10 10 
3 1 2 18 
6 1 2 3 20 18 9 
18 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
27 1 2 3 20 9 9 9 9 9 4 9 9 6 5 7 8 9 10 11 10 16 22 22 22 16 16 22 
4 1 2 18 20 
23 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 17 19 10 
3 1 2 18 
19 1 2 3 9 4 6 5 7 8 9 10 10 10 10 11 10 18 21 16 
3 1 2 18 
11 1 2 3 4 6 5 7 8 9 10 10 
6 1 2 3 9 19 9 
3 1 2 18 
4 1 2 18 20 
29 1 2 3 9 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 11 10 16 22 22 22 22 21 18 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
17 1 2 3 9 9 9 9 4 6 5 7 8 9 10 10 10 10 
17 1 2 3 20 4 5 6 7 8 9 11 10 14 15 13 12 16 
9 1 2 3 20 9 9 9 18 9 
4 1 2 18 20 
28 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 11 10 16 22 22 22 16 16 14 13 15 12 16 
13 1 2 3 9 9 9 9 9 9 9 9 19 9 
4 1 2 18 20 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
7 1 2 3 20 9 18 9 
6 1 2 3 20 19 9 
6 1 2 3 20 18 9 
3 1 2 18 
26 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 22 22 16 16 22 22 22 
10 1 2 3 20 9 9 9 9 18 9 
6 1 2 23 23 18 23 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 21 18 16 
18 1 2 3 20 4 5 6 7 8 9 10 11 10 12 13 15 14 16 
15 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
18 1 2 3 9 9 9 9 9 9 9 9 9 4 6 5 7 8 9 
34 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 22 22 22 22 22 22 22 22 22 22 22 14 15 13 12 16 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
19 1 2 3 9 9 4 5 6 7 8 9 10 11 10 14 12 15 13 16 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 14 13 15 12 16 
17 1 2 3 4 5 6 7 8 9 11 10 16 12 13 14 15 16 
6 1 2 3 20 18 9 
3 1 2 18 
5 1 2 3 18 9 
6 1 2 3 20 18 9 
8 1 2 3 9 9 9 18 9 
20 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 14 12 13 15 16 
14 1 2 3 20 4 5 6 7 8 9 10 10 10 10 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 22 13 14 12 15 16 
27 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 11 10 16 16 16 16 16 12 14 13 15 16 
3 1 2 18 
34 1 2 3 9 4 9 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 16 22 22 22 22 13 14 15 12 16 
4 1 2 18 20 
46 1 2 23 23 23 20 23 23 23 3 20 4 6 5 7 8 9 10 10 10 10 10 11 10 16 16 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 16 22 22 22 
28 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
10 1 2 3 9 9 9 9 9 19 9 
21 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 10 17 19 10 
3 1 2 18 
3 1 2 18 
14 1 2 20 3 20 9 9 9 9 9 9 9 19 9 
12 1 2 3 9 9 9 9 9 9 9 9 9 
29 1 2 3 20 9 4 5 6 7 8 9 17 5 7 8 10 11 10 16 16 22 22 22 22 13 14 12 15 16 
6 1 2 3 9 18 9 
4 1 2 18 20 
19 1 2 3 9 4 5 6 7 8 9 10 11 10 16 14 12 13 15 16 
15 1 2 3 20 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
18 1 2 3 4 5 6 7 8 9 10 10 11 10 14 13 12 15 16 
29 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 22 22 16 13 14 12 15 16 
22 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 16 
16 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 10 
4 1 2 18 20 
21 1 2 3 9 9 9 4 5 6 7 8 9 10 11 10 16 14 12 13 15 16 
21 1 2 3 20 9 9 4 6 5 7 8 9 11 10 16 23 15 13 14 12 16 
19 1 2 3 4 6 5 7 8 9 11 10 16 22 22 14 12 13 15 16 
10 1 2 3 20 9 9 9 9 18 9 
15 1 2 3 9 9 9 4 6 5 7 8 9 19 17 10 
16 1 2 3 4 6 5 7 8 9 11 10 13 14 12 15 16 
3 1 2 18 
7 1 2 3 9 9 19 9 
26 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 22 16 22 22 22 22 14 15 13 12 16 
6 1 2 3 9 19 9 
16 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 
5 1 2 3 19 9 
5 1 2 3 19 9 
6 1 2 3 9 19 9 
7 1 2 3 20 9 18 9 
15 1 2 3 20 4 6 5 7 8 9 10 10 17 19 10 
37 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 16 22 22 22 22 22 22 22 22 21 18 16 
6 1 2 3 9 19 9 
30 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 5 17 7 8 22 22 22 11 22 16 12 14 13 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
17 1 2 3 20 9 9 4 5 6 7 8 9 10 10 17 19 10 
10 1 2 3 9 9 9 9 9 18 9 
31 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
6 1 2 3 20 18 9 
5 1 2 3 18 9 
7 1 2 3 20 9 18 9 
20 1 2 3 4 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
26 1 2 3 20 9 4 5 6 7 8 9 10 10 10 11 10 16 16 16 22 22 14 12 13 15 16 
3 1 2 18 
3 1 2 18 
8 1 2 3 9 9 9 19 9 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 12 15 13 16 
17 1 2 3 9 9 4 5 6 7 8 9 10 10 10 17 19 10 
3 1 2 18 
23 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 
3 1 2 18 
5 1 2 3 18 9 
12 1 2 3 4 5 6 7 8 9 10 10 10 
19 1 2 3 20 9 9 4 6 5 7 8 9 10 10 11 10 21 18 16 
14 1 2 3 4 6 5 7 8 9 11 10 21 18 16 
3 1 2 18 
26 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 11 10 16 22 22 22 13 12 14 15 16 
33 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 16 22 22 22 16 16 13 12 14 15 16 
15 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 
20 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 13 14 12 15 16 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 11 10 16 16 12 13 15 14 16 
4 1 2 18 20 
23 1 2 3 20 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 21 18 16 
14 1 2 3 9 9 4 5 6 7 8 9 10 10 10 
18 1 2 3 9 4 5 6 7 8 9 11 10 16 14 12 13 15 16 
4 1 2 18 20 
19 1 2 3 4 5 6 7 8 9 10 10 10 11 10 14 13 12 15 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
14 1 2 20 3 20 9 9 9 9 9 9 9 9 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
13 1 2 3 9 4 5 6 7 8 9 10 10 10 
16 1 2 3 9 9 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
22 1 2 3 4 6 5 7 8 9 10 11 10 16 16 16 22 16 12 13 15 14 16 
3 1 2 18 
20 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 
13 1 2 3 9 4 5 6 7 8 9 10 10 10 
24 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 13 15 12 14 16 
12 1 2 3 4 6 5 7 8 9 19 17 10 
4 1 2 18 20 
5 1 2 3 18 9 
15 1 2 3 4 5 6 7 8 9 10 11 10 18 21 16 
22 1 2 3 9 4 6 5 7 8 9 11 10 16 16 22 22 22 22 22 18 21 16 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 19 9 
4 1 2 18 20 
6 1 2 3 20 18 9 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 13 15 12 16 
13 1 2 3 20 9 4 6 5 7 8 9 10 10 
4 1 2 18 20 
15 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 
23 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 13 14 15 12 16 
6 1 2 23 23 18 23 
16 1 2 3 9 4 5 6 7 8 9 10 11 10 21 18 16 
18 1 2 3 4 5 6 7 8 9 10 11 10 16 14 13 12 15 16 
4 1 2 18 20 
31 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 16 16 22 22 16 16 22 16 22 22 22 14 13 15 12 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 15 12 14 13 16 
3 1 2 18 
22 1 2 3 20 9 9 4 6 5 7 8 9 10 10 10 11 10 14 13 15 12 16 
5 1 2 20 18 20 
16 1 2 3 9 9 9 9 4 5 6 7 8 9 17 19 10 
3 1 2 18 
3 1 2 18 
14 1 2 3 9 9 4 5 6 7 8 9 10 10 10 
25 1 2 3 9 9 4 6 5 7 8 9 10 10 10 11 10 16 16 22 22 13 14 12 15 16 
4 1 2 18 20 
16 1 2 3 9 9 4 5 6 7 8 9 11 10 18 21 16 
21 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 16 14 12 13 15 16 
9 1 2 23 23 20 20 23 18 20 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 9 9 4 5 6 7 8 9 10 10 10 11 10 
49 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 10 10 10 11 10 16 16 16 16 16 16 16 16 22 22 22 22 22 22 22 16 22 22 22 5 17 7 8 16 22 22 22 22 22 
8 1 2 3 9 9 9 18 9 
10 1 2 3 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 4 19 9 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 10 10 10 
6 1 2 3 9 19 9 
4 1 2 18 20 
6 1 2 3 9 18 9 
6 1 2 3 4 19 9 
3 1 2 18 
24 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 16 12 14 13 15 22 
5 1 2 20 18 20 
6 1 2 3 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
15 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 
15 1 2 3 9 4 6 5 7 8 9 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
6 1 2 3 20 19 9 
30 1 2 3 20 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 16 16 16 16 16 22 22 16 21 18 16 
3 1 2 18 
28 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 16 16 16 12 13 14 15 16 
6 1 2 3 9 9 9 
28 1 2 3 9 9 9 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 16 13 14 15 12 16 
10 1 2 20 20 3 20 9 9 19 9 
3 1 2 18 
20 1 2 3 9 4 6 5 7 8 9 11 10 16 22 22 22 22 18 21 16 
17 1 2 20 3 20 9 9 4 6 5 7 8 9 10 10 10 10 
25 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 5 17 7 8 10 10 10 10 10 10 
20 1 2 3 9 4 6 5 7 8 9 17 5 7 8 10 10 10 21 18 10 
13 1 2 3 4 5 6 7 8 9 10 17 19 10 
5 1 2 20 18 20 
5 1 2 3 19 9 
3 1 2 18 
17 1 2 3 20 4 5 6 7 8 9 11 10 14 13 15 12 16 
5 1 2 3 18 9 
12 1 2 3 20 9 9 9 9 9 9 9 9 
4 1 2 18 20 
4 1 2 18 20 
12 1 2 3 9 4 5 6 7 8 9 10 10 
33 1 2 3 4 6 5 7 8 9 11 10 16 22 22 16 22 22 17 5 7 8 22 22 22 22 11 22 16 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
12 1 2 3 9 9 9 9 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
20 1 2 3 20 9 9 4 5 6 7 8 9 10 10 10 11 10 16 22 22 
7 1 2 3 20 9 18 9 
3 1 2 18 
18 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 19 9 
3 1 2 18 
17 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 
37 1 2 3 20 4 9 6 5 7 8 9 5 17 7 8 10 10 17 5 7 8 10 11 10 16 16 16 16 16 16 16 16 14 12 13 15 16 
7 1 2 3 20 9 18 9 
3 1 2 18 
14 1 2 3 20 9 9 9 9 9 9 9 9 19 9 
10 1 2 3 9 9 9 9 9 19 9 
3 1 2 18 
22 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 22 22 12 15 14 13 16 
5 1 2 3 18 9 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
15 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
23 1 2 3 4 5 6 7 8 9 10 17 5 7 8 10 10 11 10 14 12 13 15 16 
17 1 2 3 4 5 6 7 8 9 10 10 10 5 17 7 8 10 
23 1 2 3 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 
14 1 2 3 9 4 6 5 7 8 9 10 10 10 10 
6 1 2 3 20 18 9 
12 1 2 3 4 5 6 7 8 9 18 21 10 
19 1 2 3 4 6 5 7 8 9 10 11 10 16 16 22 22 21 18 22 
7 1 2 3 20 9 18 9 
3 1 2 18 
3 1 2 18 
7 1 2 3 20 9 18 9 
4 1 2 18 20 
15 1 2 3 20 9 4 5 6 7 8 9 10 10 11 10 
4 1 2 18 20 
12 1 2 3 9 4 5 6 7 8 9 10 10 
13 1 2 3 9 4 5 6 7 8 9 10 10 10 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 18 9 
7 1 2 3 9 9 18 9 
17 1 2 3 9 4 5 6 7 8 9 11 10 15 13 12 14 16 
4 1 2 18 20 
9 1 2 3 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 10 10 10 
4 1 2 18 20 
17 1 2 3 4 5 6 7 8 9 10 11 10 16 16 18 21 22 
3 1 2 18 
26 1 2 3 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 17 5 7 8 10 10 10 10 
5 1 2 3 19 9 
3 1 2 18 
5 1 2 20 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
11 1 2 3 9 9 9 9 9 9 9 9 
5 1 2 3 19 9 
14 1 2 3 4 5 6 7 8 9 10 10 17 19 10 
3 1 2 18 
4 1 2 18 20 
5 1 2 3 18 9 
13 1 2 3 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 9 9 9 9 
3 1 2 18 
40 1 2 3 9 9 9 9 9 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 11 10 16 22 22 22 22 22 22 22 14 13 12 15 16 
25 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 13 12 14 15 22 
7 1 2 3 20 9 19 9 
3 1 2 18 
12 1 2 3 4 6 5 7 8 9 17 19 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
28 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 22 22 22 22 22 22 16 22 14 12 13 15 22 
19 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 16 16 22 22 
3 1 2 18 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 13 14 12 15 16 
25 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 16 21 18 16 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 19 9 
3 1 2 18 
23 1 2 3 9 9 9 9 9 4 6 5 7 8 9 11 10 16 23 14 13 12 15 16 
27 1 2 3 4 6 5 7 8 9 5 17 7 8 10 11 10 16 17 5 7 8 16 14 13 15 12 22 
13 1 2 3 20 4 5 6 7 8 9 10 10 10 
19 1 2 3 9 9 4 5 6 7 8 9 11 10 16 22 22 21 18 16 
3 1 2 18 
23 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
22 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 11 10 16 21 18 16 
5 1 2 20 18 20 
3 1 2 18 
21 1 2 3 20 4 6 5 7 8 9 17 5 7 8 10 10 10 10 10 11 10 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
7 1 2 3 20 4 18 9 
3 1 2 18 
8 1 2 3 9 9 9 18 9 
16 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 
3 1 2 18 
22 1 2 20 3 20 9 9 4 6 5 7 8 9 10 11 10 16 13 14 15 12 16 
11 1 2 3 9 4 6 5 7 8 9 10 
21 1 2 3 4 6 5 7 8 9 11 10 16 16 22 22 22 14 12 13 15 16 
21 1 2 20 3 20 9 4 5 6 7 8 9 10 10 11 10 13 12 14 15 16 
4 1 2 18 20 
7 1 2 3 9 9 18 9 
21 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 10 10 10 10 10 
20 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 
15 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 
11 1 2 3 9 9 9 9 9 9 18 9 
3 1 2 18 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
6 1 2 3 20 19 9 
25 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 14 13 15 12 16 
3 1 2 18 
31 1 2 3 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 5 17 7 8 16 15 13 12 14 22 
3 1 2 18 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 21 18 22 
34 1 2 20 20 3 20 9 4 6 5 7 8 9 10 10 11 10 16 22 22 22 16 16 16 16 16 16 16 16 12 14 13 15 16 
6 1 2 3 20 19 9 
6 1 2 3 20 19 9 
10 1 2 3 9 9 9 9 9 19 9 
6 1 2 3 9 18 9 
25 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 
24 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 16 16 13 12 14 15 16 
3 1 2 18 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 11 10 16 22 22 14 13 12 15 16 
15 1 2 3 9 9 4 6 5 7 8 9 10 10 10 10 
10 1 2 3 9 9 9 9 4 19 9 
26 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 11 10 16 16 16 16 14 15 12 13 16 
5 1 2 20 18 20 
5 1 2 20 18 20 
6 1 2 3 9 18 9 
6 1 2 3 9 18 9 
3 1 2 18 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 13 15 12 16 
40 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 5 17 7 8 10 17 5 7 8 10 10 10 17 5 7 8 10 17 5 7 8 10 10 10 
6 1 2 3 9 19 9 
4 1 2 18 20 
17 1 2 3 4 6 5 7 8 9 11 10 16 14 13 15 12 16 
3 1 2 18 
3 1 2 18 
5 1 2 20 18 20 
23 1 2 20 3 20 9 9 9 9 4 6 5 7 8 9 10 11 10 14 12 13 15 16 
4 1 2 18 20 
20 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 13 14 12 15 16 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 
22 1 2 3 20 9 9 9 4 6 5 7 8 9 10 10 10 10 10 10 17 19 10 
13 1 2 3 9 9 9 9 9 9 9 9 9 9 
7 1 2 20 20 20 18 20 
4 1 2 18 20 
6 1 2 3 9 19 9 
3 1 2 18 
6 1 2 3 9 19 9 
14 1 2 3 20 4 5 6 7 8 9 10 10 10 10 
3 1 2 18 
15 1 2 20 3 20 9 9 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
13 1 2 3 20 4 6 5 7 8 9 10 10 10 
31 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 10 10 
4 1 2 18 20 
18 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 
17 1 2 20 20 3 20 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
11 1 2 3 9 4 5 6 7 8 9 10 
12 1 2 3 4 5 6 7 8 9 17 19 10 
3 1 2 18 
5 1 2 3 19 9 
19 1 2 20 3 20 9 4 5 6 7 8 9 10 11 10 16 18 21 16 
12 1 2 3 4 5 6 7 8 9 19 17 10 
4 1 2 18 20 
3 1 2 18 
33 1 2 3 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 16 22 22 22 16 16 16 16 15 13 14 12 16 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
14 1 2 20 20 3 20 9 9 9 9 9 9 18 9 
3 1 2 18 
3 1 2 18 
15 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 
37 1 2 3 9 4 5 6 7 8 9 10 11 10 16 16 16 16 16 22 22 22 17 5 7 8 22 22 22 22 22 11 22 15 14 13 12 16 
3 1 2 18 
13 1 2 3 9 9 4 5 6 7 8 9 10 10 
15 1 2 3 9 9 4 5 6 7 8 9 10 19 17 10 
29 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 17 5 7 8 22 22 22 22 11 22 16 
3 1 2 18 
16 1 2 3 20 9 9 9 9 9 9 9 9 9 9 19 9 
49 1 2 3 20 9 4 6 5 7 8 9 10 10 10 5 17 7 8 10 17 5 7 8 10 10 11 10 16 16 16 16 16 22 22 22 22 16 22 22 22 22 22 22 22 14 12 13 15 22 
11 1 2 3 9 9 9 9 9 9 19 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
6 1 2 3 20 18 9 
20 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 15 13 12 14 16 
31 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 16 22 22 22 22 22 22 
22 1 2 3 20 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 11 10 
22 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 16 16 14 15 12 13 16 
4 1 2 18 20 
23 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 10 11 10 
12 1 2 3 9 4 6 5 7 8 9 10 10 
21 1 2 3 20 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 
31 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 22 22 22 22 16 16 16 16 22 22 16 14 15 13 12 16 
3 1 2 18 
33 1 2 3 9 9 9 4 5 6 7 8 9 11 10 16 22 22 22 22 5 17 7 8 22 22 22 11 22 14 15 13 12 16 
18 1 2 3 9 4 5 6 7 8 9 10 10 10 11 10 18 21 16 
16 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
13 1 2 3 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
3 1 2 18 
12 1 2 3 20 9 9 9 9 9 9 9 9 
4 1 2 18 20 
3 1 2 18 
13 1 2 3 4 5 6 7 8 9 10 10 10 10 
3 1 2 18 
17 1 2 3 9 9 9 9 4 5 6 7 8 9 10 19 17 10 
30 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 17 5 7 8 10 17 5 7 8 10 10 10 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 11 10 15 13 12 14 16 
3 1 2 18 
25 1 2 3 20 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 17 5 7 8 10 10 
4 1 2 18 20 
3 1 2 18 
20 1 2 3 9 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 10 
3 1 2 18 
7 1 2 3 20 9 18 9 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 10 11 10 16 15 14 12 13 16 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
27 1 2 3 9 4 6 5 7 8 9 10 10 10 11 10 16 22 22 22 22 22 22 15 12 13 14 22 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
18 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 21 18 16 
4 1 2 18 20 
20 1 2 3 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 
3 1 2 18 
24 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 22 22 16 14 13 12 15 16 
15 1 2 3 4 5 6 7 8 9 11 10 16 18 21 16 
3 1 2 18 
3 1 2 18 
3 1 2 18 
11 1 2 3 4 6 5 7 8 9 10 10 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
21 1 2 3 9 9 9 9 4 5 6 7 8 9 10 11 10 14 13 15 12 16 
13 1 2 3 4 6 5 7 8 9 10 10 10 10 
4 1 2 18 20 
23 1 2 3 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 16 22 22 22 22 
12 1 2 3 4 5 6 7 8 9 10 10 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 9 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
6 1 2 3 9 19 9 
17 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 10 10 
4 1 2 18 20 
17 1 2 20 20 3 20 4 6 5 7 8 9 10 10 10 11 10 
5 1 2 3 18 9 
3 1 2 18 
27 1 2 3 20 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 22 22 22 12 15 13 14 16 
3 1 2 18 
17 1 2 3 9 4 5 6 7 8 9 10 10 10 10 17 19 10 
6 1 2 3 9 19 9 
3 1 2 18 
15 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 
24 1 2 20 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 10 10 10 19 17 10 
9 1 2 3 20 9 9 9 18 9 
19 1 2 3 9 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
5 1 2 3 19 9 
3 1 2 18 
21 1 2 3 9 4 6 5 7 8 9 10 5 17 7 8 10 10 10 10 10 10 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 19 17 10 
23 1 2 3 9 9 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 18 21 16 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 14 12 13 15 16 
28 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 16 16 16 22 22 19 17 22 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 9 
4 1 2 3 9 
6 1 2 20 20 18 20 
7 1 2 3 9 9 18 9 
14 1 2 3 9 9 4 6 5 7 8 9 17 19 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
20 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 11 10 18 21 16 
25 1 2 20 3 20 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 13 14 15 12 16 
5 1 2 20 18 20 
3 1 2 18 
24 1 2 3 4 5 6 7 8 9 10 11 10 16 16 5 17 7 8 16 13 14 12 15 22 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 
15 1 2 3 9 4 6 5 7 8 9 10 10 19 17 10 
14 1 2 3 9 9 4 6 5 7 8 9 10 10 10 
22 1 2 3 20 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 10 
20 1 2 3 20 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 
4 1 2 18 20 
12 1 2 3 4 5 6 7 8 9 10 10 10 
20 1 2 3 20 9 4 6 5 7 8 9 10 10 11 10 14 12 13 15 16 
3 1 2 18 
20 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 14 15 13 12 16 
16 1 2 3 20 4 6 5 7 8 9 10 10 10 10 11 10 
4 1 2 18 20 
3 1 2 18 
31 1 2 3 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 11 10 5 17 7 8 16 13 14 12 15 22 
18 1 2 3 9 9 9 9 9 9 9 4 6 5 7 8 9 10 10 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
5 1 2 20 18 20 
7 1 2 3 9 9 19 9 
17 1 2 3 4 6 5 7 8 9 10 10 17 5 7 8 10 10 
4 1 2 18 20 
22 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 22 22 16 16 17 19 16 
20 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 13 14 12 15 16 
3 1 2 18 
8 1 2 3 20 9 9 19 9 
9 1 2 3 20 9 9 9 18 9 
3 1 2 18 
20 1 2 3 4 6 5 7 8 9 10 11 10 16 16 22 22 16 16 22 22 
19 1 2 3 9 4 5 6 7 8 9 11 10 16 16 13 14 12 15 16 
3 1 2 18 
16 1 2 3 9 4 6 5 7 8 9 10 11 10 17 19 16 
14 1 2 3 20 4 6 5 7 8 9 10 10 10 10 
23 1 2 3 9 4 5 6 7 8 9 10 11 10 16 22 22 22 22 15 14 12 13 16 
5 1 2 3 18 9 
13 1 2 3 4 5 6 7 8 9 10 10 10 10 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
40 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 16 22 17 5 7 8 22 22 22 22 22 22 22 11 22 16 16 14 13 12 15 16 
7 1 2 3 9 4 19 9 
3 1 2 18 
3 1 2 18 
15 1 2 3 4 5 6 7 8 9 10 10 10 19 17 10 
3 1 2 18 
7 1 2 3 20 9 18 9 
6 1 2 3 20 18 9 
4 1 2 18 20 
4 1 2 18 20 
17 1 2 3 9 9 9 9 9 4 5 6 7 8 9 10 10 10 
3 1 2 18 
20 1 2 3 4 5 6 7 8 9 10 10 10 10 11 10 14 13 12 15 16 
17 1 2 3 4 5 6 7 8 9 10 11 10 13 12 14 15 16 
10 1 2 3 9 9 9 9 9 19 9 
7 1 2 3 20 9 19 9 
22 1 2 3 20 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 17 19 10 
13 1 2 3 4 6 5 7 8 9 10 19 17 10 
12 1 2 3 4 5 6 7 8 9 10 10 10 
3 1 2 18 
19 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 16 18 21 22 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
21 1 2 3 9 4 6 5 7 8 9 11 10 16 16 16 16 13 14 12 15 16 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
18 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 16 16 22 
22 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 11 10 15 13 12 14 16 
5 1 2 20 18 20 
5 1 2 3 18 9 
15 1 2 3 9 9 4 5 6 7 8 9 10 10 10 10 
3 1 2 18 
10 1 2 3 9 9 9 9 9 19 9 
13 1 2 3 9 4 5 6 7 8 9 10 10 10 
22 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 
3 1 2 18 
9 1 2 3 9 9 9 9 9 9 
19 1 2 3 9 9 9 9 4 5 6 7 8 9 10 11 10 21 18 16 
17 1 2 20 3 20 9 9 9 9 9 9 4 6 5 7 8 9 
39 1 2 3 9 9 4 6 5 7 8 9 17 5 7 8 10 10 11 10 16 22 22 22 16 22 22 22 22 16 17 5 7 8 16 14 15 12 13 22 
3 1 2 18 
19 1 2 3 4 6 5 7 8 9 10 5 17 7 8 10 10 19 17 10 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
7 1 2 3 9 9 19 9 
22 1 2 3 20 4 5 6 7 8 9 11 10 16 22 22 22 16 15 14 12 13 16 
15 1 2 3 20 9 4 6 5 7 8 9 10 10 10 10 
6 1 2 3 20 18 9 
3 1 2 18 
24 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 
5 1 2 20 18 20 
5 1 2 3 18 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
10 1 2 3 9 9 9 9 9 19 9 
6 1 2 3 9 9 9 
13 1 2 3 9 9 4 6 5 7 8 9 10 10 
19 1 2 3 20 9 9 9 9 9 4 6 5 7 8 9 10 10 10 10 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 14 13 12 15 16 
9 1 2 3 20 9 9 9 19 9 
20 1 2 3 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 
5 1 2 3 19 9 
26 1 2 3 4 5 6 7 8 9 11 10 16 22 22 22 22 16 16 22 22 22 14 12 13 15 16 
21 1 2 3 9 9 9 4 5 6 7 8 9 17 5 7 8 10 10 10 11 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
28 1 2 3 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 5 17 7 8 16 14 13 15 12 22 
20 1 2 3 20 9 9 9 9 4 6 5 7 8 9 10 11 10 21 18 16 
20 1 2 3 4 6 5 7 8 9 11 10 16 22 22 16 14 13 15 12 16 
18 1 2 3 20 9 9 4 6 5 7 8 9 17 5 7 8 10 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
19 1 2 3 20 9 9 9 9 9 9 4 5 6 7 8 9 10 11 10 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 20 9 9 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 
19 1 2 3 4 5 6 7 8 9 5 17 7 8 10 10 10 10 11 10 
3 1 2 18 
14 1 2 3 9 4 6 5 7 8 9 10 19 17 10 
6 1 2 3 20 18 9 
18 1 2 3 20 9 4 6 5 7 8 9 5 17 7 8 10 10 10 
3 1 2 18 
31 1 2 3 4 5 6 7 8 9 10 11 10 16 16 16 16 16 16 16 16 16 16 5 17 7 8 22 22 22 11 22 
6 1 2 3 20 18 9 
20 1 2 3 4 6 5 7 8 9 11 10 16 22 22 22 15 13 12 14 16 
12 1 2 3 9 9 9 9 9 9 9 9 9 
16 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 10 
24 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 16 16 22 22 14 12 15 13 16 
17 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
23 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 13 14 15 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
16 1 2 3 20 9 9 9 9 9 4 6 5 7 8 9 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
13 1 2 3 9 9 4 6 5 7 8 9 10 10 
3 1 2 18 
21 1 2 3 4 5 6 7 8 9 11 10 16 16 22 22 22 14 15 12 13 16 
3 1 2 18 
5 1 2 3 18 9 
3 1 2 18 
14 1 2 3 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
14 1 2 3 20 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 22 22 17 19 22 
5 1 2 20 18 20 
24 1 2 3 9 4 6 5 7 8 9 10 10 10 10 10 10 10 10 10 10 10 10 10 10 
17 1 2 3 4 5 6 7 8 9 10 11 10 16 22 17 19 22 
24 1 2 3 20 9 4 6 5 7 8 9 10 11 10 16 16 22 22 16 15 13 12 14 16 
30 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 10 11 10 17 5 7 8 16 14 13 12 15 22 
6 1 2 3 9 18 9 
16 1 2 3 9 9 9 9 9 9 9 9 9 9 4 19 9 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
16 1 2 3 9 4 6 5 7 8 9 10 17 5 7 8 10 
22 1 2 3 9 4 6 5 7 8 9 10 11 10 16 16 16 16 15 14 12 13 16 
3 1 2 18 
20 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 14 13 12 15 16 
13 1 2 3 9 9 4 6 5 7 8 9 10 10 
3 1 2 18 
13 1 2 3 4 5 6 7 8 9 10 10 11 10 
19 1 2 3 4 5 6 7 8 9 11 10 16 16 22 12 14 13 15 22 
4 1 2 18 20 
19 1 2 3 9 9 9 9 4 5 6 7 8 9 10 10 11 10 16 22 
5 1 2 3 18 9 
3 1 2 18 
15 1 2 3 20 4 6 5 7 8 9 10 10 19 17 10 
6 1 2 3 9 18 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
5 1 2 3 19 9 
4 1 2 18 20 
8 1 2 3 20 9 9 18 9 
4 1 2 18 20 
6 1 2 23 23 18 23 
11 1 2 3 9 4 5 6 7 8 9 10 
17 1 2 3 9 4 6 5 7 8 9 11 10 14 12 13 15 16 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 13 12 14 15 16 
19 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 10 10 10 
18 1 2 3 9 4 5 6 7 8 9 10 11 10 13 14 15 12 16 
3 1 2 18 
6 1 2 3 9 18 9 
38 1 2 3 9 9 4 6 5 7 8 9 10 10 11 10 16 16 22 22 22 22 22 22 22 22 22 22 22 16 22 22 22 22 22 22 22 22 22 
15 1 2 3 4 6 5 7 8 9 10 11 10 21 18 16 
4 1 2 18 20 
6 1 2 3 20 19 9 
3 1 2 18 
7 1 2 3 9 9 19 9 
40 1 2 3 9 9 9 4 6 5 7 8 9 17 5 7 8 10 10 10 5 17 7 8 10 17 5 7 8 10 10 10 17 5 7 8 10 10 10 11 10 
18 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 11 10 
28 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 11 10 5 17 7 8 16 13 14 15 12 22 
3 1 2 18 
9 1 2 3 9 9 9 9 19 9 
9 1 2 3 9 9 9 9 19 9 
10 1 2 3 9 9 9 9 9 18 9 
12 1 2 3 9 4 5 6 7 8 9 10 10 
7 1 2 3 9 9 19 9 
3 1 2 18 
37 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 17 5 7 8 10 17 5 7 8 10 11 10 16 22 22 14 15 12 13 16 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 14 12 15 16 
17 1 2 3 20 9 9 9 9 4 5 6 7 8 9 10 10 10 
10 1 2 3 4 9 9 9 9 9 9 
3 1 2 18 
19 1 2 3 20 9 9 9 9 4 6 5 7 8 9 11 10 18 21 16 
21 1 2 3 4 6 5 7 8 9 10 10 10 11 10 16 16 16 22 22 22 22 
11 1 2 3 4 6 5 7 8 9 10 10 
22 1 2 3 9 9 4 6 5 7 8 9 5 17 7 8 10 10 10 10 10 10 10 
4 1 2 18 20 
29 1 2 3 9 9 9 9 4 6 5 7 8 9 11 10 16 16 16 16 16 16 5 17 7 8 22 22 22 22 
21 1 2 3 20 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 
12 1 2 3 9 4 6 5 7 8 9 10 10 
3 1 2 18 
26 1 2 3 9 9 4 6 5 7 8 9 10 11 10 16 22 22 22 22 22 16 14 15 12 13 16 
12 1 2 3 20 4 6 5 7 8 9 10 10 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
9 1 2 3 20 9 9 9 18 9 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
8 1 2 3 20 9 9 18 9 
3 1 2 18 
3 1 2 18 
15 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 
3 1 2 18 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 10 10 10 
22 1 2 3 4 5 6 7 8 9 11 10 16 16 16 22 22 22 14 12 13 15 16 
3 1 2 18 
18 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 19 9 
3 1 2 18 
36 1 2 3 20 4 5 6 7 8 9 10 10 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 22 14 13 12 15 22 
3 1 2 18 
3 1 2 18 
3 1 2 18 
16 1 2 3 4 5 6 7 8 9 17 5 7 8 10 10 10 
10 1 2 20 3 20 9 9 9 18 9 
5 1 2 3 18 9 
12 1 2 3 20 4 6 5 7 8 9 10 10 
9 1 2 3 20 9 9 9 18 9 
17 1 2 3 9 9 9 4 6 5 7 8 9 10 10 10 11 10 
27 1 2 3 4 6 5 7 8 9 10 10 10 10 5 17 7 8 10 11 10 16 16 14 15 12 13 16 
3 1 2 18 
12 1 2 3 9 4 6 5 7 8 9 10 10 
20 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
4 1 2 18 20 
11 1 2 3 4 5 6 7 8 9 10 10 
14 1 2 3 20 4 6 5 7 8 9 10 11 10 16 
3 1 2 18 
20 1 2 3 20 4 5 6 7 8 9 10 11 10 16 16 12 13 15 14 16 
13 1 2 3 4 6 5 7 8 9 10 10 11 10 
47 1 2 3 9 9 9 9 9 9 4 9 9 5 6 7 8 9 5 17 7 8 10 10 11 10 16 22 5 17 7 8 22 22 22 22 22 22 22 22 22 11 22 15 13 12 14 16 
21 1 2 3 9 9 9 4 5 6 7 8 9 10 17 5 7 8 10 10 11 10 
17 1 2 3 4 6 5 7 8 9 10 11 10 12 13 15 14 16 
8 1 2 3 9 9 9 9 9 
8 1 2 3 9 9 9 18 9 
53 1 2 3 9 9 9 9 9 4 5 6 7 8 9 17 5 7 8 10 5 17 7 8 10 5 17 7 8 10 10 10 10 17 5 7 8 10 10 11 10 5 17 7 8 16 11 22 16 15 12 14 13 22 
3 1 2 18 
15 1 2 3 9 9 9 4 5 6 7 8 9 10 10 10 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
17 1 2 3 4 5 6 7 8 9 10 11 10 12 13 15 14 16 
3 1 2 18 
14 1 2 3 9 4 6 5 7 8 9 10 10 11 10 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 12 13 15 16 
4 1 2 18 20 
19 1 2 3 9 9 4 6 5 7 8 9 11 10 16 15 12 13 14 16 
17 1 2 3 4 5 6 7 8 9 10 11 10 14 13 12 15 16 
3 1 2 18 
16 1 2 3 9 9 9 9 9 4 6 5 7 8 9 10 10 
18 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
3 1 2 18 
3 1 2 18 
7 1 2 3 9 9 19 9 
13 1 2 3 20 9 9 9 9 9 9 9 9 9 
15 1 2 3 4 6 5 7 8 9 10 11 10 21 18 16 
23 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
26 1 2 3 9 4 6 5 7 8 9 11 10 16 17 5 7 8 22 22 11 22 14 12 15 13 16 
4 1 2 18 20 
14 1 2 3 20 9 4 5 6 7 8 9 10 11 10 
6 1 2 3 20 18 9 
18 1 2 3 9 4 6 5 7 8 9 10 11 10 12 14 13 15 16 
3 1 2 18 
13 1 2 3 20 9 9 9 9 9 9 9 18 9 
6 1 2 23 23 18 23 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
5 1 2 3 20 9 
3 1 2 18 
3 1 2 18 
16 1 2 3 4 6 5 7 8 9 17 5 7 8 10 10 10 
8 1 2 3 20 9 9 18 9 
5 1 2 3 18 9 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
6 1 2 20 20 18 20 
12 1 2 3 4 5 6 7 8 9 10 10 10 
17 1 2 20 3 20 9 9 9 4 5 6 7 8 9 10 10 10 
4 1 2 18 20 
3 1 2 18 
18 1 2 3 20 9 4 5 6 7 8 9 11 10 13 12 14 15 16 
17 1 2 3 9 4 5 6 7 8 9 11 10 14 15 13 12 16 
7 1 2 3 20 9 18 9 
3 1 2 18 
44 1 2 3 9 9 9 4 6 5 7 8 9 10 11 10 16 16 16 16 22 22 16 16 16 16 16 22 22 22 5 17 7 8 22 22 11 22 16 16 12 13 15 14 16 
4 1 2 18 20 
25 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 17 5 7 8 10 10 11 10 
3 1 2 18 
11 1 2 3 4 5 6 7 8 9 10 10 
30 1 2 3 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 16 16 16 16 22 22 22 13 14 12 15 16 
3 1 2 18 
17 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 
5 1 2 3 18 9 
14 1 2 3 9 9 9 9 9 9 9 9 9 19 9 
13 1 2 3 9 9 9 4 5 6 7 8 9 10 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
12 1 2 3 4 5 6 7 8 9 10 10 10 
3 1 2 18 
3 1 2 18 
21 1 2 3 9 9 4 5 6 7 8 9 10 10 11 10 16 16 22 22 22 22 
4 1 2 18 20 
4 1 2 18 20 
11 1 2 3 4 5 6 7 8 9 10 10 
22 1 2 3 9 9 4 5 6 7 8 9 11 10 16 16 22 22 12 13 15 14 22 
21 1 2 3 9 9 9 9 4 6 5 7 8 9 10 11 10 14 12 13 15 16 
4 1 2 18 20 
4 1 2 18 20 
10 1 2 3 20 9 9 9 9 18 9 
3 1 2 18 
21 1 2 20 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
20 1 2 3 4 6 5 7 8 9 10 10 11 10 16 16 13 14 12 15 16 
16 1 2 3 9 4 5 6 7 8 9 10 10 10 10 11 10 
13 1 2 3 9 9 4 5 6 7 8 9 10 10 
5 1 2 20 18 20 
14 1 2 3 9 4 5 6 7 8 9 10 17 19 10 
7 1 2 3 20 9 18 9 
24 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 22 22 22 22 16 22 21 18 22 
12 1 2 3 4 6 5 7 8 9 10 10 10 
3 1 2 18 
23 1 2 3 20 4 6 5 7 8 9 10 10 11 10 16 16 16 16 15 13 14 12 16 
3 1 2 18 
13 1 2 3 9 4 5 6 7 8 9 19 17 10 
13 1 2 3 9 4 5 6 7 8 9 10 11 10 
3 1 2 18 
6 1 2 3 9 18 9 
47 1 2 3 20 4 6 5 7 8 9 10 11 10 17 5 7 8 16 22 22 22 22 22 22 22 22 11 22 16 16 22 16 22 22 22 22 22 22 17 5 7 8 22 22 22 22 22 
5 1 2 20 18 20 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 18 9 
4 1 2 18 20 
12 1 2 3 4 6 5 7 8 9 10 10 10 
7 1 2 3 9 9 19 9 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
16 1 2 3 4 5 6 7 8 9 11 10 16 16 18 21 16 
16 1 2 3 20 9 9 4 6 5 7 8 9 10 10 11 10 
13 1 2 3 9 4 5 6 7 8 9 10 11 10 
3 1 2 18 
3 1 2 18 
3 1 2 18 
37 1 2 3 20 9 9 4 5 6 7 8 9 10 11 10 16 16 22 22 22 22 22 22 22 22 22 16 16 16 16 16 17 5 7 8 22 22 
12 1 2 3 20 9 9 9 9 9 9 18 9 
20 1 2 3 9 4 6 5 7 8 9 10 11 10 16 22 13 12 14 15 22 
17 1 2 3 9 4 5 6 7 8 9 10 10 11 10 21 18 16 
13 1 2 20 20 3 20 9 9 9 9 9 9 9 
4 1 2 18 20 
4 1 2 18 20 
20 1 2 3 20 9 9 9 4 5 6 7 8 9 11 10 16 16 21 18 16 
12 1 2 3 4 6 5 7 8 9 10 11 10 
3 1 2 18 
11 1 2 3 20 4 6 5 7 8 9 10 
3 1 2 18 
6 1 2 3 9 18 9 
27 1 2 3 20 4 5 6 7 8 9 17 5 7 8 10 10 11 10 16 16 16 16 13 14 12 15 16 
23 1 2 3 4 5 6 7 8 9 10 11 10 16 22 22 22 16 16 14 13 15 12 16 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 11 10 
8 1 2 20 3 20 9 19 9 
4 1 2 18 20 
17 1 2 23 20 23 23 23 23 23 23 20 3 20 9 9 18 9 
12 1 2 3 4 5 6 7 8 9 10 10 10 
3 1 2 18 
23 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 
11 1 2 3 9 4 6 5 7 8 9 10 
8 1 2 3 9 9 9 19 9 
3 1 2 18 
6 1 2 20 20 18 20 
21 1 2 3 20 9 9 9 9 9 9 9 9 9 9 4 5 6 7 8 9 10 
18 1 2 3 4 6 5 7 8 9 10 11 10 16 14 12 13 15 16 
4 1 2 18 20 
14 1 2 3 20 9 9 4 6 5 7 8 9 10 10 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 9 9 4 5 6 7 8 9 5 17 7 8 10 10 
14 1 2 3 4 5 6 7 8 9 10 11 10 16 22 
17 1 2 3 9 9 9 9 9 9 9 9 4 5 6 7 8 9 
3 1 2 18 
21 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 11 10 21 18 16 
3 1 2 18 
19 1 2 3 9 4 5 6 7 8 9 10 11 10 16 14 15 13 12 22 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
13 1 2 3 4 6 5 7 8 9 10 10 11 10 
6 1 2 20 20 18 20 
14 1 2 20 3 20 9 9 4 5 6 7 8 9 10 
20 1 2 3 9 4 5 6 7 8 9 11 10 16 22 22 14 12 13 15 16 
3 1 2 18 
7 1 2 3 20 9 18 9 
11 1 2 3 9 4 6 5 7 8 9 10 
15 1 2 20 3 20 9 4 5 6 7 8 9 10 10 10 
4 1 2 18 20 
14 1 2 3 20 9 9 4 6 5 7 8 9 11 10 
4 1 2 18 20 
15 1 2 3 20 4 5 6 7 8 9 11 10 18 21 16 
16 1 2 3 20 9 9 4 6 5 7 8 9 10 10 11 10 
19 1 2 3 9 4 5 6 7 8 9 10 17 5 7 8 10 10 11 10 
13 1 2 3 9 4 6 5 7 8 9 10 11 10 
11 1 2 3 4 6 5 7 8 9 10 10 
13 1 2 3 9 9 9 9 9 9 9 9 9 9 
8 1 2 3 9 9 9 19 9 
16 1 2 3 9 9 9 9 9 9 4 5 6 7 8 9 10 
7 1 2 3 20 9 18 9 
8 1 2 3 9 9 9 19 9 
3 1 2 18 
4 1 2 18 20 
22 1 2 3 20 4 6 5 7 8 9 10 11 10 16 16 22 22 14 12 13 15 16 
17 1 2 3 9 9 9 4 5 6 7 8 9 5 17 7 8 10 
7 1 2 3 9 9 9 9 
11 1 2 20 3 20 9 9 9 9 18 9 
3 1 2 18 
19 1 2 3 9 4 5 6 7 8 9 11 10 16 16 14 15 12 13 16 
3 1 2 18 
3 1 2 18 
21 1 2 3 20 9 9 9 4 5 6 7 8 9 10 11 10 14 13 15 12 16 
20 1 2 3 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 10 10 
24 1 2 3 9 4 6 5 7 8 9 10 10 10 10 11 10 16 22 22 22 22 21 18 22 
11 1 2 3 9 4 5 6 7 8 9 10 
20 1 2 20 3 20 9 4 5 6 7 8 9 5 17 7 8 10 10 10 10 
13 1 2 3 4 5 6 7 8 9 10 19 17 10 
12 1 2 3 4 5 6 7 8 9 19 17 10 
22 1 2 3 9 9 4 5 6 7 8 9 10 11 10 16 16 16 13 12 14 15 16 
3 1 2 18 
36 1 2 3 20 4 6 5 7 8 9 11 10 16 22 22 22 22 22 22 22 22 22 22 22 22 22 16 16 22 22 22 22 22 22 16 22 
3 1 2 18 
22 1 2 3 9 9 4 6 5 7 8 9 11 10 16 22 22 22 14 12 13 15 16 
13 1 2 3 9 9 9 4 5 6 7 8 9 10 
20 1 2 3 20 9 9 4 6 5 7 8 9 10 11 10 14 13 12 15 16 
25 1 2 3 20 4 5 6 7 8 9 10 17 5 7 8 10 10 10 11 10 16 16 21 18 16 
10 1 2 3 4 6 5 7 8 9 10 
4 1 2 18 20 
11 1 2 3 4 6 5 7 8 9 10 10 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
3 1 2 18 
17 1 2 3 20 4 6 5 7 8 9 11 10 13 14 12 15 16 
14 1 2 3 4 5 6 7 8 9 10 10 10 10 10 
17 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 16 22 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
12 1 2 3 9 9 4 5 6 7 8 9 10 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
17 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
5 1 2 20 18 20 
8 1 2 3 20 9 9 18 9 
6 1 2 3 20 18 9 
6 1 2 3 20 18 9 
4 1 2 18 20 
31 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 11 10 16 16 22 22 22 22 22 22 14 15 12 13 16 
15 1 2 3 9 4 5 6 7 8 9 11 10 21 18 16 
3 1 2 18 
14 1 2 3 4 5 6 7 8 9 10 10 19 17 10 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
3 1 2 18 
26 1 2 3 4 6 5 7 8 9 11 10 16 17 5 7 8 16 22 22 22 22 22 22 22 22 22 
19 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
3 1 2 18 
25 1 2 3 20 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
23 1 2 3 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 19 9 
4 1 2 18 20 
13 1 2 3 20 9 9 4 6 5 7 8 9 10 
25 1 2 3 9 4 5 6 7 8 9 17 5 7 8 10 10 10 17 5 7 8 10 10 11 10 
12 1 2 3 4 5 6 7 8 9 10 10 10 
3 1 2 18 
3 1 2 18 
19 1 2 3 4 5 6 7 8 9 10 11 10 16 23 13 14 12 15 16 
14 1 2 3 9 9 9 4 5 6 7 8 9 10 10 
24 1 2 3 9 9 4 5 6 7 8 9 11 10 16 22 22 22 16 16 14 13 12 15 16 
3 1 2 18 
4 1 2 18 20 
6 1 2 20 20 18 20 
20 1 2 3 9 4 5 6 7 8 9 10 10 11 10 16 15 13 12 14 16 
17 1 2 3 4 6 5 7 8 9 10 17 5 7 8 10 10 10 
9 1 2 3 20 9 9 9 18 9 
17 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 
17 1 2 3 4 6 5 7 8 9 10 11 10 13 12 14 15 16 
3 1 2 18 
5 1 2 3 19 9 
4 1 2 18 20 
10 1 2 3 4 5 6 7 8 9 10 
4 1 2 18 20 
23 1 2 3 9 9 9 4 6 5 7 8 9 11 10 16 16 22 16 12 15 14 13 16 
10 1 2 3 9 9 9 9 9 19 9 
5 1 2 3 18 9 
19 1 2 3 9 4 5 6 7 8 9 10 11 10 16 14 15 13 12 16 
3 1 2 18 
13 1 2 3 9 4 5 6 7 8 9 10 10 10 
24 1 2 3 9 4 5 6 7 8 9 11 10 16 16 5 17 7 8 16 22 22 22 22 22 
18 1 2 3 4 5 6 7 8 9 10 5 17 7 8 10 10 10 10 
3 1 2 18 
3 1 2 18 
6 1 2 3 9 19 9 
5 1 2 20 18 20 
9 1 2 3 9 9 9 9 9 9 
3 1 2 18 
12 1 2 3 9 9 4 6 5 7 8 9 10 
17 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 
3 1 2 18 
6 1 2 3 20 18 9 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
3 1 2 18 
4 1 2 18 20 
4 1 2 18 20 
3 1 2 18 
4 1 2 18 20 
9 1 2 3 9 9 9 9 9 9 
4 1 2 18 20 
13 1 2 3 4 5 6 7 8 9 10 11 10 16 
14 1 2 3 9 9 9 4 6 5 7 8 9 11 10 
11 1 2 3 9 4 5 6 7 8 9 10 
18 1 2 3 9 4 6 5 7 8 9 10 10 11 10 16 18 21 16 
19 1 2 3 9 4 6 5 7 8 9 5 17 7 8 10 10 10 11 10 
3 1 2 18 
4 1 2 18 20 
11 1 2 3 20 4 5 6 7 8 9 10 
4 1 2 18 20 
