1434 28
4 1 2 3 2 
9 1 4 2 3 2 5 3 2 3 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 8 9 10 11 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 5 7 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
10 1 2 6 7 4 16 17 18 4 5 
1 1 
6 1 2 6 7 4 5 
7 1 2 6 7 4 5 12 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 4 5 7 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
5 1 2 6 7 4 
1 1 
4 1 2 4 6 
6 1 2 6 4 5 7 
1 1 
1 1 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
1 1 
6 1 2 6 7 4 5 
1 1 
1 1 
5 1 2 6 4 7 
1 1 
1 1 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
3 1 4 16 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
10 1 2 6 7 4 5 12 13 14 15 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 8 9 10 11 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 8 9 10 11 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
5 1 2 6 7 4 
4 1 2 6 7 
4 1 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
4 1 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
3 1 4 5 
6 1 2 6 7 4 5 
5 1 2 6 7 4 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
4 1 2 6 7 
6 1 2 6 7 4 5 
6 1 4 2 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 4 5 8 9 10 11 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 4 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
10 1 2 6 4 5 8 9 10 11 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 4 2 6 7 5 8 9 10 11 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
4 1 2 6 7 
4 1 2 6 7 
4 1 2 6 7 
8 1 4 2 16 4 5 6 7 
8 1 4 5 2 3 2 6 7 
14 1 4 2 3 2 19 4 5 3 2 3 2 6 7 
10 1 4 2 6 7 17 19 20 4 5 
6 1 2 4 5 6 7 
10 1 2 4 5 3 2 3 2 6 7 
6 1 2 6 7 4 5 
8 1 4 21 4 5 2 6 7 
8 1 2 3 2 6 4 5 7 
14 1 4 19 16 17 18 21 22 23 2 6 7 4 5 
6 1 4 5 2 6 7 
9 1 4 5 12 13 2 6 7 24 
6 1 2 6 7 4 5 
6 1 4 2 6 5 7 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
8 1 4 5 2 3 2 6 7 
1 1 
6 1 2 6 7 4 5 
10 1 4 5 2 3 2 3 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
1 1 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
10 1 4 5 8 9 10 11 2 6 7 
1 1 
8 1 4 5 2 3 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
8 1 4 5 2 3 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
8 1 2 3 2 6 7 4 5 
6 1 4 5 2 6 7 
10 1 2 4 3 2 3 2 6 7 19 
1 1 
12 1 4 19 4 5 2 3 2 3 2 6 7 
6 1 4 5 2 6 7 
8 1 2 3 2 6 7 4 5 
6 1 4 5 2 6 7 
8 1 2 4 16 4 6 7 5 
6 1 2 6 7 4 5 
8 1 4 5 2 3 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
8 1 2 3 2 6 7 4 5 
6 1 4 5 2 6 7 
10 1 4 4 4 22 4 5 2 6 7 
6 1 2 4 6 5 7 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
5 1 2 6 3 4 
10 1 4 19 4 19 4 5 2 6 7 
13 1 4 5 2 3 2 3 2 6 3 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
9 1 4 17 20 4 5 2 6 7 
1 1 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 4 2 5 6 7 
6 1 4 5 2 6 7 
1 1 
6 1 4 2 5 6 7 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 4 6 7 5 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
8 1 2 6 7 4 16 4 5 
1 1 
1 1 
1 1 
1 1 
1 1 
6 1 2 6 4 5 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
1 1 
1 1 
6 1 4 2 6 7 5 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 4 5 7 
6 1 2 6 4 7 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
12 1 4 5 12 13 2 6 7 24 13 14 15 
6 1 2 4 5 6 7 
10 1 2 6 4 5 7 12 13 14 15 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
12 1 2 6 4 19 4 19 4 19 4 5 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
12 1 2 6 7 4 19 4 5 8 9 10 11 
6 1 2 4 5 6 7 
10 1 4 16 17 18 4 5 2 6 7 
6 1 4 2 6 7 5 
6 1 2 4 5 6 7 
9 1 2 6 7 4 16 22 4 5 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 4 2 5 6 7 
5 1 2 6 7 4 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 4 2 6 5 7 
12 1 4 5 8 9 10 11 2 3 2 6 7 
6 1 2 6 7 4 5 
5 1 2 6 7 4 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 4 5 7 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
10 1 4 5 2 6 7 12 13 14 15 
6 1 4 5 2 6 7 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 5 6 7 
6 1 2 6 4 5 7 
6 1 4 2 6 5 7 
6 1 2 4 6 5 7 
6 1 2 6 7 4 5 
10 1 2 6 7 4 19 4 19 4 5 
6 1 2 6 4 5 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
12 1 4 23 17 25 4 23 4 5 2 6 7 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
15 1 2 6 7 4 21 23 4 21 23 4 21 23 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
18 1 2 6 4 7 23 4 23 4 23 4 23 4 23 4 23 4 5 
6 1 2 6 4 5 7 
6 1 2 6 4 7 5 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
7 1 2 6 4 5 7 12 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
8 1 2 6 4 16 4 5 7 
8 1 4 5 2 3 2 6 7 
8 1 2 6 7 4 16 4 5 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
8 1 4 23 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
18 1 2 6 4 19 4 19 4 19 4 19 4 7 19 4 19 4 5 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
9 1 4 2 6 17 18 4 5 7 
6 1 2 4 5 6 7 
6 1 4 2 5 6 7 
6 1 4 5 2 6 7 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 4 6 5 7 
6 1 2 4 6 7 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
5 1 2 6 7 4 
6 1 2 6 7 4 5 
1 1 
12 1 2 6 4 23 7 4 23 4 23 4 5 
6 1 2 6 7 4 5 
8 1 2 4 16 4 5 6 7 
6 1 4 5 2 6 7 
12 1 4 23 4 23 2 6 4 23 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
1 1 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
1 1 
6 1 2 6 7 4 5 
10 1 2 4 16 4 16 4 5 6 7 
6 1 4 5 2 6 7 
12 1 4 5 2 3 2 3 2 3 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 2 6 4 5 7 
1 1 
6 1 4 5 2 6 7 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
8 1 4 19 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
8 1 4 5 2 3 2 6 7 
1 1 
10 1 2 6 7 4 16 4 16 4 5 
6 1 2 4 6 7 5 
6 1 4 5 2 6 7 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
1 1 
8 1 4 16 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
1 1 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
12 1 2 4 16 4 16 4 16 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
1 1 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
1 1 
5 1 4 5 2 6 
7 1 4 5 2 6 7 12 
1 1 
1 1 
1 1 
1 1 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
1 1 
6 1 2 4 5 6 7 
10 1 2 6 7 4 5 8 9 10 11 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 4 5 7 
10 1 2 4 5 12 13 6 14 7 15 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
1 1 
1 1 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
11 1 4 2 6 7 17 20 4 16 4 5 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
8 1 2 4 16 4 5 6 7 
1 1 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
1 1 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
1 1 
8 1 4 16 23 4 16 2 23 
6 1 2 6 7 4 5 
13 1 4 17 16 23 18 4 5 2 3 2 6 7 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
8 1 2 3 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
10 1 2 6 4 16 4 16 4 5 7 
6 1 2 4 6 5 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 5 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 4 7 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
1 1 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
10 1 2 6 4 5 8 9 10 11 7 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 4 16 4 16 4 5 6 7 
6 1 2 6 7 4 5 
8 1 4 16 4 5 2 6 7 
6 1 2 6 7 4 5 
8 1 2 6 4 16 4 5 7 
9 1 4 23 16 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 4 6 7 5 12 13 14 15 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
1 1 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
1 1 
6 1 4 2 5 6 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
5 1 2 6 7 4 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
10 1 2 4 5 6 7 12 13 14 15 
10 1 2 6 7 4 5 12 13 14 15 
5 1 2 6 7 4 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
18 1 2 6 7 4 5 8 9 26 9 26 9 26 9 26 9 10 11 
6 1 4 2 6 7 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 4 2 6 7 5 
6 1 2 4 5 6 7 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
9 1 2 6 7 4 17 18 4 5 
6 1 4 5 2 6 7 
6 1 2 4 6 7 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 4 6 5 7 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 8 9 10 11 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
3 1 4 2 
8 1 2 4 19 4 5 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 2 4 6 7 5 
6 1 2 6 4 5 7 
1 1 
6 1 2 4 5 6 7 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
7 1 2 6 4 5 7 12 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 4 2 6 7 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
8 1 4 5 2 3 2 6 7 
1 1 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
4 1 2 4 3 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 4 5 2 6 7 
6 1 2 6 4 5 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
9 1 4 19 16 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
1 1 
1 1 
6 1 2 6 7 4 5 
1 1 
12 1 2 6 7 4 19 4 19 4 19 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
5 1 2 6 7 4 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 4 2 5 6 7 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 4 2 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 16 17 20 4 5 
1 1 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 4 2 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 4 6 7 5 
8 1 2 6 7 4 23 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 8 9 10 11 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 4 6 5 7 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
6 1 2 4 6 5 7 
6 1 2 4 5 6 7 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 4 2 6 7 5 12 13 14 15 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
8 1 4 2 6 7 23 4 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 4 5 7 
6 1 2 4 5 6 7 
6 1 2 6 4 7 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 4 5 2 6 7 12 13 14 15 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
10 1 4 5 2 6 7 8 9 10 11 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 4 5 6 7 
1 1 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 4 6 7 5 
6 1 2 6 4 7 5 
6 1 2 4 6 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
14 1 2 6 7 4 5 8 9 26 9 26 9 10 11 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
6 1 2 6 4 5 7 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
5 1 2 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
16 1 2 3 2 3 2 3 2 3 2 3 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
8 1 2 3 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 4 5 7 
10 1 2 4 4 4 5 3 2 6 7 
6 1 2 6 4 5 7 
1 1 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
7 1 2 4 5 6 3 2 
18 1 2 6 7 4 17 25 18 21 19 27 20 23 16 22 4 4 4 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
4 1 2 3 2 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 4 7 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 4 2 6 7 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
3 1 2 4 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
9 1 2 4 6 3 2 5 6 7 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
24 1 4 2 16 6 7 4 16 4 16 4 16 4 16 4 16 4 16 4 16 4 16 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 4 5 7 
6 1 2 4 5 6 7 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 7 5 
3 1 4 2 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
8 1 2 3 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
3 1 2 4 
6 1 2 6 7 4 5 
1 1 
1 1 
1 1 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 4 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 5 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
5 1 2 6 7 4 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
18 1 2 3 2 3 2 6 7 4 16 4 16 4 5 12 13 14 15 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
1 1 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
5 1 2 6 7 4 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
12 1 2 6 7 4 21 23 4 23 21 4 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 4 6 7 19 17 25 4 5 
6 1 2 6 7 4 5 
3 1 4 2 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 3 2 3 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 4 5 2 6 7 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 5 7 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
5 1 2 6 7 4 
25 1 2 4 17 25 6 3 2 6 7 23 4 17 25 23 4 23 17 25 4 17 25 23 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
10 1 2 4 5 12 6 7 13 14 15 
10 1 2 4 5 6 7 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
9 1 2 6 7 4 17 25 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 8 9 10 11 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 4 5 6 7 12 13 14 15 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 8 9 10 11 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 4 5 2 6 7 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 5 2 6 7 
1 1 
6 1 4 5 2 6 7 
6 1 2 6 7 4 5 
10 1 4 2 6 5 7 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
6 1 2 6 4 7 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 12 13 14 15 
10 1 2 6 7 4 5 12 13 14 15 
6 1 2 4 6 5 7 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 4 2 5 6 7 
1 1 
1 1 
6 1 2 6 7 4 5 
1 1 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
4 1 4 5 2 
1 1 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
1 1 
3 1 4 2 
8 1 4 22 4 5 2 6 7 
1 1 
6 1 2 6 4 5 7 
6 1 2 6 7 4 5 
8 1 2 6 7 4 22 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
10 1 2 6 4 7 5 12 13 14 15 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 5 6 7 
10 1 2 6 7 4 5 8 9 10 11 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 2 4 5 6 7 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 4 6 7 5 
6 1 2 6 7 4 5 
10 1 2 6 7 4 5 8 9 10 11 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
9 1 2 4 5 6 3 2 6 7 
6 1 4 2 6 7 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
6 1 2 6 7 4 5 
